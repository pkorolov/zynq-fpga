module Control(input clk, input reset,
    output[2:0] io_dpath_sel_pc,
    output io_dpath_killd,
    output io_dpath_ren_1,
    output io_dpath_ren_0,
    output[2:0] io_dpath_sel_alu2,
    output[1:0] io_dpath_sel_alu1,
    output[2:0] io_dpath_sel_imm,
    output io_dpath_fn_dw,
    output[3:0] io_dpath_fn_alu,
    output io_dpath_div_mul_val,
    output io_dpath_div_mul_kill,
    //output io_dpath_div_val
    //output io_dpath_div_kill
    output[2:0] io_dpath_csr,
    output io_dpath_sret,
    output io_dpath_mem_load,
    output io_dpath_wb_load,
    output io_dpath_ex_fp_val,
    output io_dpath_mem_fp_val,
    output io_dpath_ex_wen,
    output io_dpath_ex_valid,
    output io_dpath_mem_jalr,
    output io_dpath_mem_branch,
    output io_dpath_mem_wen,
    output io_dpath_wb_wen,
    output[2:0] io_dpath_ex_mem_type,
    output io_dpath_ex_rs2_val,
    output io_dpath_ex_rocc_val,
    output io_dpath_mem_rocc_val,
    output io_dpath_bypass_1,
    output io_dpath_bypass_0,
    output[1:0] io_dpath_bypass_src_1,
    output[1:0] io_dpath_bypass_src_0,
    output io_dpath_ll_ready,
    output io_dpath_retire,
    output io_dpath_exception,
    output[63:0] io_dpath_cause,
    output io_dpath_badvaddr_wen,
    input [31:0] io_dpath_inst,
    //input  io_dpath_jalr_eq
    input  io_dpath_mem_br_taken,
    input  io_dpath_mem_misprediction,
    input  io_dpath_div_mul_rdy,
    input  io_dpath_ll_wen,
    input [4:0] io_dpath_ll_waddr,
    input [4:0] io_dpath_ex_waddr,
    input  io_dpath_mem_rs1_ra,
    input [4:0] io_dpath_mem_waddr,
    input [4:0] io_dpath_wb_waddr,
    input [7:0] io_dpath_status_ip,
    input [7:0] io_dpath_status_im,
    input [6:0] io_dpath_status_zero,
    input  io_dpath_status_er,
    input  io_dpath_status_vm,
    input  io_dpath_status_s64,
    input  io_dpath_status_u64,
    input  io_dpath_status_ef,
    input  io_dpath_status_pei,
    input  io_dpath_status_ei,
    input  io_dpath_status_ps,
    input  io_dpath_status_s,
    input  io_dpath_fp_sboard_clr,
    input [4:0] io_dpath_fp_sboard_clra,
    input  io_dpath_csr_replay,
    output io_imem_req_valid,
    //output[43:0] io_imem_req_bits_pc
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input [42:0] io_imem_btb_resp_bits_target,
    input [2:0] io_imem_btb_resp_bits_entry,
    input [3:0] io_imem_btb_resp_bits_bht_index,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output[42:0] io_imem_btb_update_bits_prediction_bits_target,
    output[2:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[3:0] io_imem_btb_update_bits_prediction_bits_bht_index,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    //output[42:0] io_imem_btb_update_bits_pc
    //output[42:0] io_imem_btb_update_bits_target
    //output[42:0] io_imem_btb_update_bits_returnAddr
    output io_imem_btb_update_bits_taken,
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isCall,
    output io_imem_btb_update_bits_isReturn,
    output io_imem_btb_update_bits_incorrectTarget,
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    output io_imem_invalidate,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output io_dmem_req_bits_kill,
    output[2:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_phys,
    //output[43:0] io_dmem_req_bits_addr
    //output[63:0] io_dmem_req_bits_data
    //output[7:0] io_dmem_req_bits_tag
    output[4:0] io_dmem_req_bits_cmd,
    input  io_dmem_resp_valid,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [2:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [7:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    //output io_dtlb_val
    //output io_dtlb_kill
    //input  io_dtlb_rdy
    //input  io_dtlb_miss
    //input  io_xcpt_dtlb_ld
    //input  io_xcpt_dtlb_st
    output io_fpu_valid,
    //input  io_fpu_fcsr_rdy
    input  io_fpu_nack_mem,
    input  io_fpu_illegal_rm,
    output io_fpu_killx,
    output io_fpu_killm,
    //input [4:0] io_fpu_dec_cmd
    //input  io_fpu_dec_ldst
    input  io_fpu_dec_wen,
    input  io_fpu_dec_ren1,
    input  io_fpu_dec_ren2,
    input  io_fpu_dec_ren3,
    //input  io_fpu_dec_swap23
    //input  io_fpu_dec_single
    //input  io_fpu_dec_fromint
    //input  io_fpu_dec_toint
    //input  io_fpu_dec_fastpipe
    //input  io_fpu_dec_fma
    //input  io_fpu_dec_round
    //input  io_fpu_sboard_set
    //input  io_fpu_sboard_clr
    //input [4:0] io_fpu_sboard_clra
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[3:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [3:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    output io_rocc_exception
);

  wire T0;
  reg  wb_reg_xcpt;
  wire T1;
  wire T2;
  wire take_pc_wb;
  wire T3;
  reg  wb_reg_sret;
  wire T4;
  wire T5;
  wire T6;
  reg  mem_reg_replay;
  wire T7;
  wire replay_ex;
  wire replay_ex_other;
  reg  mem_reg_replay_next;
  wire T8;
  reg  ex_reg_replay_next;
  wire T9;
  wire T10;
  wire id_csr_flush;
  wire T11;
  wire T12;
  wire T13;
  wire[11:0] T14;
  wire[11:0] T15;
  wire T16;
  wire[11:0] T17;
  wire T18;
  wire id_csr_wen;
  wire T19;
  wire T20;
  wire T21;
  wire[1:0] T22;
  wire T23;
  wire[31:0] T24;
  wire T25;
  wire[31:0] T26;
  wire T27;
  wire T28;
  wire[4:0] T29;
  wire T30;
  wire T31;
  wire[31:0] T32;
  wire ctrl_killd;
  wire T33;
  wire ctrl_draind;
  wire id_interrupt;
  wire id_interrupt_unmasked;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire ctrl_stalld;
  wire id_do_fence;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[31:0] T70;
  wire T71;
  wire T72;
  wire[31:0] T73;
  wire T74;
  wire T75;
  wire[31:0] T76;
  wire T77;
  wire T78;
  wire[31:0] T79;
  wire T80;
  wire T81;
  wire[31:0] T82;
  wire T83;
  wire[31:0] T84;
  reg  id_reg_fence;
  wire T85;
  wire T86;
  wire T87;
  wire id_mem_busy;
  reg  ex_reg_mem_val;
  wire T88;
  wire T89;
  wire T90;
  wire id_fence_next;
  wire T91;
  wire T92;
  wire T93;
  wire[31:0] T94;
  wire T95;
  wire[31:0] T96;
  wire T97;
  wire T98;
  wire[31:0] T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire id_sboard_hazard;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire[4:0] T110;
  wire[4:0] T111;
  wire[4:0] T112;
  wire T113;
  wire[31:0] T114;
  wire[31:0] T115;
  wire[31:0] T116;
  wire[31:0] T117;
  reg [31:0] R118;
  wire[31:0] T119;
  wire[31:0] T120;
  wire[31:0] T121;
  wire[31:0] T122;
  wire[31:0] T123;
  wire[31:0] T124;
  wire T125;
  wire wb_set_sboard;
  reg  wb_reg_rocc_val;
  wire T126;
  reg  mem_reg_rocc_val;
  wire T127;
  reg  ex_reg_rocc_val;
  wire T128;
  wire T129;
  wire ctrl_killx;
  wire T130;
  wire take_pc_mem_wb;
  wire take_pc_mem;
  wire T131;
  reg  mem_reg_jal;
  wire T132;
  reg  ex_reg_jal;
  wire T133;
  wire T134;
  wire[31:0] T135;
  wire T136;
  reg  mem_reg_jalr;
  wire T137;
  reg  ex_reg_jalr;
  wire T138;
  wire T139;
  wire[31:0] T140;
  reg  mem_reg_branch;
  wire T141;
  reg  ex_reg_branch;
  wire T142;
  wire T143;
  wire[31:0] T144;
  wire ctrl_killm;
  wire T145;
  wire fpu_kill_mem;
  reg  mem_reg_fp_val;
  wire T146;
  reg  ex_reg_fp_val;
  wire T147;
  wire T148;
  wire mem_xcpt;
  wire T149;
  reg  mem_reg_mem_val;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  reg  mem_reg_xcpt;
  wire T158;
  wire ex_xcpt;
  wire T159;
  wire T160;
  reg  ex_reg_xcpt;
  wire T161;
  wire id_xcpt;
  wire T162;
  wire[31:0] T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire[31:0] T168;
  wire T169;
  wire id_csr_privileged;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire[1:0] T175;
  wire T176;
  wire T177;
  wire[1:0] T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire[1:0] T183;
  wire T184;
  wire T185;
  wire[1:0] T186;
  wire T187;
  wire T188;
  wire[1:0] T189;
  wire T190;
  wire T191;
  wire id_csr_invalid;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire[31:0] T273;
  wire T274;
  wire T275;
  wire[31:0] T276;
  wire T277;
  wire T278;
  wire[31:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[31:0] T284;
  wire T285;
  wire T286;
  wire[31:0] T287;
  wire T288;
  wire T289;
  wire[31:0] T290;
  wire T291;
  wire T292;
  wire[31:0] T293;
  wire T294;
  wire T295;
  wire[31:0] T296;
  wire T297;
  wire T298;
  wire T299;
  wire[31:0] T300;
  wire T301;
  wire T302;
  wire[31:0] T303;
  wire T304;
  wire T305;
  wire[31:0] T306;
  wire T307;
  wire T308;
  wire[31:0] T309;
  wire T310;
  wire T311;
  wire[31:0] T312;
  wire T313;
  wire T314;
  wire[31:0] T315;
  wire T316;
  wire T317;
  wire[31:0] T318;
  wire T319;
  wire T320;
  wire[31:0] T321;
  wire T322;
  wire T323;
  wire[31:0] T324;
  wire T325;
  wire T326;
  wire[31:0] T327;
  wire T328;
  wire T329;
  wire[31:0] T330;
  wire T331;
  wire T332;
  wire[31:0] T333;
  wire T334;
  wire T335;
  wire T336;
  reg  ex_reg_xcpt_interrupt;
  wire T337;
  wire T338;
  wire T339;
  reg  mem_reg_xcpt_interrupt;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire killm_common;
  wire T344;
  reg  mem_reg_valid;
  wire T345;
  reg  ex_reg_valid;
  wire T346;
  wire T347;
  wire T348;
  wire dcache_kill_mem;
  reg  mem_reg_wen;
  wire T349;
  reg  ex_reg_wen;
  wire T350;
  wire T351;
  wire T352;
  wire[31:0] T353;
  wire T354;
  wire T355;
  wire[31:0] T356;
  wire T357;
  wire T358;
  wire[31:0] T359;
  wire T360;
  wire T361;
  wire[31:0] T362;
  wire T363;
  wire T364;
  wire T365;
  wire[31:0] T366;
  wire T367;
  wire[31:0] T368;
  wire T369;
  wire wb_dcache_miss;
  wire T370;
  reg  wb_reg_mem_val;
  wire T371;
  reg  wb_reg_div_mul_val;
  wire T372;
  reg  mem_reg_div_mul_val;
  wire T373;
  reg  ex_reg_div_mul_val;
  wire T374;
  wire T375;
  wire T376;
  wire[31:0] T377;
  wire T378;
  wire[31:0] T379;
  wire T380;
  wire id_wen_not0;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire[4:0] T387;
  wire[4:0] T388;
  wire[4:0] T389;
  wire T390;
  wire id_renx2_not0;
  wire T391;
  wire T392;
  wire T393;
  wire[31:0] T394;
  wire T395;
  wire T396;
  wire[31:0] T397;
  wire T398;
  wire[31:0] T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire[4:0] T404;
  wire[4:0] T405;
  wire T406;
  wire id_renx1_not0;
  wire T407;
  wire T408;
  wire T409;
  wire[31:0] T410;
  wire T411;
  wire T412;
  wire[31:0] T413;
  wire T414;
  wire T415;
  wire[31:0] T416;
  wire T417;
  wire T418;
  wire[31:0] T419;
  wire T420;
  wire[31:0] T421;
  wire T422;
  wire id_wb_hazard;
  wire T423;
  wire T424;
  reg  wb_reg_fp_val;
  wire T425;
  wire fp_data_hazard_wb;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire[4:0] T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  reg  wb_reg_fp_wen;
  wire T438;
  reg  mem_reg_fp_wen;
  wire T439;
  reg  ex_reg_fp_wen;
  wire T440;
  wire T441;
  wire data_hazard_wb;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  reg  wb_reg_wen;
  wire T450;
  wire T451;
  wire id_mem_hazard;
  wire T452;
  wire fp_data_hazard_mem;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  reg  mem_reg_slow_bypass;
  wire T470;
  wire ex_slow_bypass;
  wire T471;
  wire T472;
  reg [2:0] ex_reg_mem_type;
  wire[2:0] T473;
  wire[2:0] T474;
  wire[2:0] T475;
  wire[1:0] T476;
  wire T477;
  wire[31:0] T478;
  wire T479;
  wire[31:0] T480;
  wire T481;
  wire[31:0] T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  reg [4:0] ex_reg_mem_cmd;
  wire[4:0] T490;
  wire[4:0] T491;
  wire[3:0] T492;
  wire[2:0] T493;
  wire[1:0] T494;
  wire T495;
  wire T496;
  wire[31:0] T497;
  wire T498;
  wire T499;
  wire[31:0] T500;
  wire T501;
  wire[31:0] T502;
  wire T503;
  wire T504;
  wire[31:0] T505;
  wire T506;
  wire[31:0] T507;
  wire T508;
  wire T509;
  wire[31:0] T510;
  wire T511;
  wire T512;
  wire[31:0] T513;
  wire T514;
  wire[31:0] T515;
  wire T516;
  wire T517;
  reg [1:0] mem_reg_csr;
  wire[1:0] T518;
  reg [1:0] ex_reg_csr;
  wire[1:0] T519;
  wire data_hazard_mem;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire id_ex_hazard;
  wire T528;
  wire T529;
  wire fp_data_hazard_ex;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire data_hazard_ex;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  reg  ex_reg_load_use;
  wire T559;
  wire id_load_use;
  wire T560;
  wire T561;
  wire replay_ex_structural;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  reg  mem_reg_sret;
  wire T567;
  reg  ex_reg_sret;
  wire T568;
  wire T569;
  wire replay_wb;
  wire T570;
  wire T571;
  wire replay_wb_common;
  wire T572;
  reg  wb_reg_replay;
  wire T573;
  wire T574;
  wire replay_mem;
  wire T575;
  wire wb_rocc_val;
  wire T576;
  wire T577;
  reg  wb_reg_flush_inst;
  wire T578;
  reg  mem_reg_flush_inst;
  wire T579;
  reg  ex_reg_flush_inst;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  reg [1:0] mem_reg_btb_resp_bht_value;
  wire[1:0] T587;
  reg [1:0] ex_reg_btb_resp_bht_value;
  wire[1:0] T588;
  wire T589;
  wire T590;
  reg  ex_reg_btb_hit;
  wire T591;
  reg [3:0] mem_reg_btb_resp_bht_index;
  wire[3:0] T592;
  reg [3:0] ex_reg_btb_resp_bht_index;
  wire[3:0] T593;
  reg [2:0] mem_reg_btb_resp_entry;
  wire[2:0] T594;
  reg [2:0] ex_reg_btb_resp_entry;
  wire[2:0] T595;
  reg [42:0] mem_reg_btb_resp_target;
  wire[42:0] T596;
  reg [42:0] ex_reg_btb_resp_target;
  wire[42:0] T597;
  reg  mem_reg_btb_resp_taken;
  wire T598;
  reg  ex_reg_btb_resp_taken;
  wire T599;
  reg  mem_reg_btb_hit;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  reg [63:0] wb_reg_cause;
  wire[63:0] T605;
  wire[63:0] mem_cause;
  wire[63:0] T606;
  wire[3:0] T607;
  wire[3:0] T608;
  wire[3:0] T609;
  reg [63:0] mem_reg_cause;
  wire[63:0] T610;
  wire[63:0] ex_cause;
  reg [63:0] ex_reg_cause;
  wire[63:0] T611;
  wire[63:0] id_cause;
  wire[63:0] T612;
  wire[3:0] T613;
  wire[3:0] T614;
  wire[3:0] T615;
  wire[3:0] T616;
  wire[3:0] T617;
  wire[3:0] T618;
  wire[63:0] id_interrupt_cause;
  wire[63:0] T619;
  wire[63:0] T620;
  wire[63:0] T621;
  wire[63:0] T622;
  wire[63:0] T623;
  wire[63:0] T624;
  wire T625;
  wire T626;
  reg  wb_reg_valid;
  wire T627;
  wire T628;
  wire[1:0] T629;
  wire[1:0] T630;
  wire[1:0] T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire[1:0] T639;
  wire[1:0] T640;
  wire[1:0] T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire[2:0] T670;
  reg [1:0] wb_reg_csr;
  wire[1:0] T671;
  wire T672;
  wire[3:0] T673;
  wire[3:0] T674;
  wire[2:0] T675;
  wire[1:0] T676;
  wire T677;
  wire T678;
  wire[31:0] T679;
  wire T680;
  wire T681;
  wire[31:0] T682;
  wire T683;
  wire[31:0] T684;
  wire T685;
  wire T686;
  wire[31:0] T687;
  wire T688;
  wire T689;
  wire[31:0] T690;
  wire T691;
  wire T692;
  wire[31:0] T693;
  wire T694;
  wire T695;
  wire[31:0] T696;
  wire T697;
  wire[31:0] T698;
  wire T699;
  wire T700;
  wire[31:0] T701;
  wire T702;
  wire T703;
  wire[31:0] T704;
  wire T705;
  wire T706;
  wire[31:0] T707;
  wire T708;
  wire[31:0] T709;
  wire T710;
  wire T711;
  wire[31:0] T712;
  wire T713;
  wire T714;
  wire T715;
  wire[31:0] T716;
  wire T717;
  wire T718;
  wire T719;
  wire[31:0] T720;
  wire T721;
  wire[31:0] T722;
  wire[2:0] T723;
  wire[2:0] T724;
  wire[1:0] T725;
  wire T726;
  wire T727;
  wire[31:0] T728;
  wire T729;
  wire[31:0] T730;
  wire T731;
  wire T732;
  wire[31:0] T733;
  wire T734;
  wire T735;
  wire[31:0] T736;
  wire T737;
  wire T738;
  wire[31:0] T739;
  wire[1:0] T740;
  wire[1:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire[31:0] T746;
  wire T747;
  wire[31:0] T748;
  wire T749;
  wire T750;
  wire[31:0] T751;
  wire[2:0] T752;
  wire[1:0] T753;
  wire[1:0] T754;
  wire T755;
  wire T756;
  wire[31:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire T761;
  wire[31:0] T762;
  wire T763;
  wire[31:0] T764;
  wire T765;
  wire T766;
  wire[31:0] T767;
  wire T768;
  wire T769;
  wire T770;
  wire[31:0] T771;
  wire T772;
  wire T773;
  wire T774;
  wire[2:0] T775;
  wire[1:0] T776;
  wire[1:0] T777;
  wire[1:0] T778;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    wb_reg_xcpt = {1{$random}};
    wb_reg_sret = {1{$random}};
    mem_reg_replay = {1{$random}};
    mem_reg_replay_next = {1{$random}};
    ex_reg_replay_next = {1{$random}};
    id_reg_fence = {1{$random}};
    ex_reg_mem_val = {1{$random}};
    R118 = {1{$random}};
    wb_reg_rocc_val = {1{$random}};
    mem_reg_rocc_val = {1{$random}};
    ex_reg_rocc_val = {1{$random}};
    mem_reg_jal = {1{$random}};
    ex_reg_jal = {1{$random}};
    mem_reg_jalr = {1{$random}};
    ex_reg_jalr = {1{$random}};
    mem_reg_branch = {1{$random}};
    ex_reg_branch = {1{$random}};
    mem_reg_fp_val = {1{$random}};
    ex_reg_fp_val = {1{$random}};
    mem_reg_mem_val = {1{$random}};
    mem_reg_xcpt = {1{$random}};
    ex_reg_xcpt = {1{$random}};
    ex_reg_xcpt_interrupt = {1{$random}};
    mem_reg_xcpt_interrupt = {1{$random}};
    mem_reg_valid = {1{$random}};
    ex_reg_valid = {1{$random}};
    mem_reg_wen = {1{$random}};
    ex_reg_wen = {1{$random}};
    wb_reg_mem_val = {1{$random}};
    wb_reg_div_mul_val = {1{$random}};
    mem_reg_div_mul_val = {1{$random}};
    ex_reg_div_mul_val = {1{$random}};
    wb_reg_fp_val = {1{$random}};
    wb_reg_fp_wen = {1{$random}};
    mem_reg_fp_wen = {1{$random}};
    ex_reg_fp_wen = {1{$random}};
    wb_reg_wen = {1{$random}};
    mem_reg_slow_bypass = {1{$random}};
    ex_reg_mem_type = {1{$random}};
    ex_reg_mem_cmd = {1{$random}};
    mem_reg_csr = {1{$random}};
    ex_reg_csr = {1{$random}};
    ex_reg_load_use = {1{$random}};
    mem_reg_sret = {1{$random}};
    ex_reg_sret = {1{$random}};
    wb_reg_replay = {1{$random}};
    wb_reg_flush_inst = {1{$random}};
    mem_reg_flush_inst = {1{$random}};
    ex_reg_flush_inst = {1{$random}};
    mem_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_hit = {1{$random}};
    mem_reg_btb_resp_bht_index = {1{$random}};
    ex_reg_btb_resp_bht_index = {1{$random}};
    mem_reg_btb_resp_entry = {1{$random}};
    ex_reg_btb_resp_entry = {1{$random}};
    mem_reg_btb_resp_target = {2{$random}};
    ex_reg_btb_resp_target = {2{$random}};
    mem_reg_btb_resp_taken = {1{$random}};
    ex_reg_btb_resp_taken = {1{$random}};
    mem_reg_btb_hit = {1{$random}};
    wb_reg_cause = {2{$random}};
    mem_reg_cause = {2{$random}};
    ex_reg_cause = {2{$random}};
    wb_reg_valid = {1{$random}};
    wb_reg_csr = {1{$random}};
  end
`endif

  assign io_rocc_exception = T0;
  assign T0 = wb_reg_xcpt & io_dpath_status_er;
  assign T1 = mem_xcpt & T2;
  assign T2 = take_pc_wb ^ 1'h1;
  assign take_pc_wb = T3;
  assign T3 = T569 | wb_reg_sret;
  assign T4 = ctrl_killm ? 1'h0 : T5;
  assign T5 = mem_reg_sret & T6;
  assign T6 = mem_reg_replay ^ 1'h1;
  assign T7 = T566 & replay_ex;
  assign replay_ex = replay_ex_structural | replay_ex_other;
  assign replay_ex_other = T558 | mem_reg_replay_next;
  assign T8 = ctrl_killx ? 1'h0 : ex_reg_replay_next;
  assign T9 = ctrl_killd ? 1'h0 : T10;
  assign T10 = T31 | id_csr_flush;
  assign id_csr_flush = T18 & T11;
  assign T11 = T12 ^ 1'h1;
  assign T12 = T16 | T13;
  assign T13 = T14 == 12'h0;
  assign T14 = T15 & 12'h88d;
  assign T15 = io_dpath_inst[5'h1f:5'h14];
  assign T16 = T17 == 12'h0;
  assign T17 = T15 & 12'h88e;
  assign T18 = T30 & id_csr_wen;
  assign id_csr_wen = T28 | T19;
  assign T19 = T20 ^ 1'h1;
  assign T20 = T27 | T21;
  assign T21 = 2'h3 == T22;
  assign T22 = {T25, T23};
  assign T23 = T24 == 32'h1050;
  assign T24 = io_dpath_inst & 32'h1050;
  assign T25 = T26 == 32'h2050;
  assign T26 = io_dpath_inst & 32'h2050;
  assign T27 = 2'h2 == T22;
  assign T28 = T29 != 5'h0;
  assign T29 = io_dpath_inst[5'h13:4'hf];
  assign T30 = T22 != 2'h0;
  assign T31 = T32 == 32'h1008;
  assign T32 = io_dpath_inst & 32'h3058;
  assign ctrl_killd = T33;
  assign T33 = T64 | ctrl_draind;
  assign ctrl_draind = id_interrupt | ex_reg_replay_next;
  assign id_interrupt = io_dpath_status_ei & id_interrupt_unmasked;
  assign id_interrupt_unmasked = T37 | T34;
  assign T34 = T36 & T35;
  assign T35 = io_dpath_status_ip[3'h7:3'h7];
  assign T36 = io_dpath_status_im[3'h7:3'h7];
  assign T37 = T41 | T38;
  assign T38 = T40 & T39;
  assign T39 = io_dpath_status_ip[3'h6:3'h6];
  assign T40 = io_dpath_status_im[3'h6:3'h6];
  assign T41 = T45 | T42;
  assign T42 = T44 & T43;
  assign T43 = io_dpath_status_ip[3'h5:3'h5];
  assign T44 = io_dpath_status_im[3'h5:3'h5];
  assign T45 = T49 | T46;
  assign T46 = T48 & T47;
  assign T47 = io_dpath_status_ip[3'h4:3'h4];
  assign T48 = io_dpath_status_im[3'h4:3'h4];
  assign T49 = T53 | T50;
  assign T50 = T52 & T51;
  assign T51 = io_dpath_status_ip[2'h3:2'h3];
  assign T52 = io_dpath_status_im[2'h3:2'h3];
  assign T53 = T57 | T54;
  assign T54 = T56 & T55;
  assign T55 = io_dpath_status_ip[2'h2:2'h2];
  assign T56 = io_dpath_status_im[2'h2:2'h2];
  assign T57 = T61 | T58;
  assign T58 = T60 & T59;
  assign T59 = io_dpath_status_ip[1'h1:1'h1];
  assign T60 = io_dpath_status_im[1'h1:1'h1];
  assign T61 = T63 & T62;
  assign T62 = io_dpath_status_ip[1'h0:1'h0];
  assign T63 = io_dpath_status_im[1'h0:1'h0];
  assign T64 = T556 | ctrl_stalld;
  assign ctrl_stalld = T102 | id_do_fence;
  assign id_do_fence = id_mem_busy & T65;
  assign T65 = T66 | id_csr_flush;
  assign T66 = T97 | T67;
  assign T67 = id_reg_fence & T68;
  assign T68 = T71 | T69;
  assign T69 = T70 == 32'h1000202f;
  assign T70 = io_dpath_inst & 32'hf9f0607f;
  assign T71 = T74 | T72;
  assign T72 = T73 == 32'h800202f;
  assign T73 = io_dpath_inst & 32'he800607f;
  assign T74 = T77 | T75;
  assign T75 = T76 == 32'h202f;
  assign T76 = io_dpath_inst & 32'h1800607f;
  assign T77 = T80 | T78;
  assign T78 = T79 == 32'h3;
  assign T79 = io_dpath_inst & 32'h107f;
  assign T80 = T83 | T81;
  assign T81 = T82 == 32'h3;
  assign T82 = io_dpath_inst & 32'h207f;
  assign T83 = T84 == 32'h3;
  assign T84 = io_dpath_inst & 32'h405f;
  assign T85 = reset ? 1'h0 : T86;
  assign T86 = id_fence_next | T87;
  assign T87 = id_reg_fence & id_mem_busy;
  assign id_mem_busy = T90 | ex_reg_mem_val;
  assign T88 = ctrl_killd ? 1'h0 : T89;
  assign T89 = T68;
  assign T90 = io_dmem_ordered ^ 1'h1;
  assign id_fence_next = T95 | T91;
  assign T91 = T93 & T92;
  assign T92 = io_dpath_inst[5'h19:5'h19];
  assign T93 = T94 == 32'h2008;
  assign T94 = io_dpath_inst & 32'h6048;
  assign T95 = T96 == 32'h8;
  assign T96 = io_dpath_inst & 32'h3058;
  assign T97 = T100 | T98;
  assign T98 = T99 == 32'h100f;
  assign T99 = io_dpath_inst & 32'h707f;
  assign T100 = T93 & T101;
  assign T101 = io_dpath_inst[5'h1a:5'h1a];
  assign T102 = T105 | T103;
  assign T103 = T68 & T104;
  assign T104 = io_dmem_req_ready ^ 1'h1;
  assign T105 = T422 | id_sboard_hazard;
  assign id_sboard_hazard = T382 | T106;
  assign T106 = id_wen_not0 & T107;
  assign T107 = T113 & T108;
  assign T108 = T109 - 1'h1;
  assign T109 = 1'h1 << T110;
  assign T110 = T111 + 5'h1;
  assign T111 = T112 - T112;
  assign T112 = io_dpath_inst[4'hb:3'h7];
  assign T113 = T114 >> T112;
  assign T114 = R118 & T115;
  assign T115 = ~ T116;
  assign T116 = io_dpath_ll_wen ? T117 : 32'h0;
  assign T117 = 1'h1 << io_dpath_ll_waddr;
  assign T119 = reset ? 32'h0 : T120;
  assign T120 = T380 ? T122 : T121;
  assign T121 = io_dpath_ll_wen ? T114 : R118;
  assign T122 = T114 | T123;
  assign T123 = T125 ? T124 : 32'h0;
  assign T124 = 1'h1 << io_dpath_wb_waddr;
  assign T125 = wb_set_sboard & io_dpath_wb_wen;
  assign wb_set_sboard = T369 | wb_reg_rocc_val;
  assign T126 = ctrl_killm ? 1'h0 : mem_reg_rocc_val;
  assign T127 = ctrl_killx ? 1'h0 : ex_reg_rocc_val;
  assign T128 = ctrl_killd ? 1'h0 : T129;
  assign T129 = 1'h0;
  assign ctrl_killx = T130;
  assign T130 = take_pc_mem_wb | replay_ex;
  assign take_pc_mem_wb = take_pc_wb | take_pc_mem;
  assign take_pc_mem = io_dpath_mem_misprediction & T131;
  assign T131 = T136 | mem_reg_jal;
  assign T132 = ctrl_killx ? 1'h0 : ex_reg_jal;
  assign T133 = ctrl_killd ? 1'h0 : T134;
  assign T134 = T135 == 32'h48;
  assign T135 = io_dpath_inst & 32'h48;
  assign T136 = mem_reg_branch | mem_reg_jalr;
  assign T137 = ctrl_killx ? 1'h0 : ex_reg_jalr;
  assign T138 = ctrl_killd ? 1'h0 : T139;
  assign T139 = T140 == 32'h4;
  assign T140 = io_dpath_inst & 32'h1c;
  assign T141 = ctrl_killx ? 1'h0 : ex_reg_branch;
  assign T142 = ctrl_killd ? 1'h0 : T143;
  assign T143 = T144 == 32'h40;
  assign T144 = io_dpath_inst & 32'h54;
  assign ctrl_killm = T145;
  assign T145 = T148 | fpu_kill_mem;
  assign fpu_kill_mem = mem_reg_fp_val & io_fpu_nack_mem;
  assign T146 = ctrl_killx ? 1'h0 : ex_reg_fp_val;
  assign T147 = ctrl_killd ? 1'h0 : 1'h0;
  assign T148 = killm_common | mem_xcpt;
  assign mem_xcpt = T151 | T149;
  assign T149 = mem_reg_mem_val & io_dmem_xcpt_pf_st;
  assign T150 = ctrl_killx ? 1'h0 : ex_reg_mem_val;
  assign T151 = T153 | T152;
  assign T152 = mem_reg_mem_val & io_dmem_xcpt_pf_ld;
  assign T153 = T155 | T154;
  assign T154 = mem_reg_mem_val & io_dmem_xcpt_ma_st;
  assign T155 = T157 | T156;
  assign T156 = mem_reg_mem_val & io_dmem_xcpt_ma_ld;
  assign T157 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign T158 = ctrl_killx ? 1'h0 : ex_xcpt;
  assign ex_xcpt = T160 | T159;
  assign T159 = ex_reg_fp_val & io_fpu_illegal_rm;
  assign T160 = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign T161 = ctrl_killd ? 1'h0 : id_xcpt;
  assign id_xcpt = T164 | T162;
  assign T162 = T163 == 32'h50;
  assign T163 = io_dpath_inst & 32'h80003050;
  assign T164 = T169 | T165;
  assign T165 = T167 & T166;
  assign T166 = io_dpath_status_s ^ 1'h1;
  assign T167 = T168 == 32'h80000050;
  assign T168 = io_dpath_inst & 32'h80003050;
  assign T169 = T190 | id_csr_privileged;
  assign id_csr_privileged = T30 & T170;
  assign T170 = T176 | T171;
  assign T171 = T172 & id_csr_wen;
  assign T172 = T174 & T173;
  assign T173 = io_dpath_status_s ^ 1'h1;
  assign T174 = T175 == 2'h1;
  assign T175 = T15[4'h9:4'h8];
  assign T176 = T179 | T177;
  assign T177 = 2'h2 <= T178;
  assign T178 = T15[4'h9:4'h8];
  assign T179 = T184 | T180;
  assign T180 = T182 & T181;
  assign T181 = io_dpath_status_s ^ 1'h1;
  assign T182 = T183 == 2'h1;
  assign T183 = T15[4'hb:4'ha];
  assign T184 = T187 | T185;
  assign T185 = T186 == 2'h2;
  assign T186 = T15[4'hb:4'ha];
  assign T187 = T188 & id_csr_wen;
  assign T188 = T189 == 2'h3;
  assign T189 = T15[4'hb:4'ha];
  assign T190 = T335 | T191;
  assign T191 = T270 | id_csr_invalid;
  assign id_csr_invalid = T30 & T192;
  assign T192 = T193 ^ 1'h1;
  assign T193 = T195 | T194;
  assign T194 = 12'hccf == T15;
  assign T195 = T197 | T196;
  assign T196 = 12'hcce == T15;
  assign T197 = T199 | T198;
  assign T198 = 12'hccd == T15;
  assign T199 = T201 | T200;
  assign T200 = 12'hccc == T15;
  assign T201 = T203 | T202;
  assign T202 = 12'hccb == T15;
  assign T203 = T205 | T204;
  assign T204 = 12'hcca == T15;
  assign T205 = T207 | T206;
  assign T206 = 12'hcc9 == T15;
  assign T207 = T209 | T208;
  assign T208 = 12'hcc8 == T15;
  assign T209 = T211 | T210;
  assign T210 = 12'hcc7 == T15;
  assign T211 = T213 | T212;
  assign T212 = 12'hcc6 == T15;
  assign T213 = T215 | T214;
  assign T214 = 12'hcc5 == T15;
  assign T215 = T217 | T216;
  assign T216 = 12'hcc4 == T15;
  assign T217 = T219 | T218;
  assign T218 = 12'hcc3 == T15;
  assign T219 = T221 | T220;
  assign T220 = 12'hcc2 == T15;
  assign T221 = T223 | T222;
  assign T222 = 12'hcc1 == T15;
  assign T223 = T225 | T224;
  assign T224 = 12'hcc0 == T15;
  assign T225 = T227 | T226;
  assign T226 = 12'hc02 == T15;
  assign T227 = T229 | T228;
  assign T228 = 12'hc01 == T15;
  assign T229 = T231 | T230;
  assign T230 = 12'hc00 == T15;
  assign T231 = T233 | T232;
  assign T232 = 12'h51f == T15;
  assign T233 = T235 | T234;
  assign T234 = 12'h51e == T15;
  assign T235 = T237 | T236;
  assign T236 = 12'h51d == T15;
  assign T237 = T239 | T238;
  assign T238 = 12'h50f == T15;
  assign T239 = T241 | T240;
  assign T240 = 12'h50e == T15;
  assign T241 = T243 | T242;
  assign T242 = 12'h50d == T15;
  assign T243 = T245 | T244;
  assign T244 = 12'h50c == T15;
  assign T245 = T247 | T246;
  assign T246 = 12'h50b == T15;
  assign T247 = T249 | T248;
  assign T248 = 12'h50a == T15;
  assign T249 = T251 | T250;
  assign T250 = 12'h509 == T15;
  assign T251 = T253 | T252;
  assign T252 = 12'h508 == T15;
  assign T253 = T255 | T254;
  assign T254 = 12'h507 == T15;
  assign T255 = T257 | T256;
  assign T256 = 12'h506 == T15;
  assign T257 = T259 | T258;
  assign T258 = 12'h505 == T15;
  assign T259 = T261 | T260;
  assign T260 = 12'h504 == T15;
  assign T261 = T263 | T262;
  assign T262 = 12'h503 == T15;
  assign T263 = T265 | T264;
  assign T264 = 12'h502 == T15;
  assign T265 = T267 | T266;
  assign T266 = 12'h501 == T15;
  assign T267 = T269 | T268;
  assign T268 = 12'h500 == T15;
  assign T269 = 12'hc0 == T15;
  assign T270 = T271 ^ 1'h1;
  assign T271 = T274 | T272;
  assign T272 = T273 == 32'h33;
  assign T273 = io_dpath_inst & 32'hfc007077;
  assign T274 = T277 | T275;
  assign T275 = T276 == 32'h4063;
  assign T276 = io_dpath_inst & 32'h407f;
  assign T277 = T280 | T278;
  assign T278 = T279 == 32'h1063;
  assign T279 = io_dpath_inst & 32'h306f;
  assign T280 = T281 | T69;
  assign T281 = T282 | T72;
  assign T282 = T285 | T283;
  assign T283 = T284 == 32'h2004033;
  assign T284 = io_dpath_inst & 32'hfe004077;
  assign T285 = T288 | T286;
  assign T286 = T287 == 32'h5033;
  assign T287 = io_dpath_inst & 32'hbe007077;
  assign T288 = T291 | T289;
  assign T289 = T290 == 32'h501b;
  assign T290 = io_dpath_inst & 32'hbe00705f;
  assign T291 = T294 | T292;
  assign T292 = T293 == 32'h5013;
  assign T293 = io_dpath_inst & 32'hbc00707f;
  assign T294 = T297 | T295;
  assign T295 = T296 == 32'h2073;
  assign T296 = io_dpath_inst & 32'h207f;
  assign T297 = T298 | T75;
  assign T298 = T301 | T299;
  assign T299 = T300 == 32'h2013;
  assign T300 = io_dpath_inst & 32'h207f;
  assign T301 = T304 | T302;
  assign T302 = T303 == 32'h101b;
  assign T303 = io_dpath_inst & 32'hfe00305f;
  assign T304 = T307 | T305;
  assign T305 = T306 == 32'h1013;
  assign T306 = io_dpath_inst & 32'hfc00305f;
  assign T307 = T310 | T308;
  assign T308 = T309 == 32'h73;
  assign T309 = io_dpath_inst & 32'h7fffffff;
  assign T310 = T313 | T311;
  assign T311 = T312 == 32'h6f;
  assign T312 = io_dpath_inst & 32'h7f;
  assign T313 = T316 | T314;
  assign T314 = T315 == 32'h63;
  assign T315 = io_dpath_inst & 32'h707b;
  assign T316 = T319 | T317;
  assign T317 = T318 == 32'h33;
  assign T318 = io_dpath_inst & 32'hbe007077;
  assign T319 = T322 | T320;
  assign T320 = T321 == 32'h33;
  assign T321 = io_dpath_inst & 32'hfc00007f;
  assign T322 = T325 | T323;
  assign T323 = T324 == 32'h17;
  assign T324 = io_dpath_inst & 32'h5f;
  assign T325 = T328 | T326;
  assign T326 = T327 == 32'h13;
  assign T327 = io_dpath_inst & 32'h7077;
  assign T328 = T331 | T329;
  assign T329 = T330 == 32'hf;
  assign T330 = io_dpath_inst & 32'h607f;
  assign T331 = T334 | T332;
  assign T332 = T333 == 32'h3;
  assign T333 = io_dpath_inst & 32'h106f;
  assign T334 = T83 | T81;
  assign T335 = T336 | io_imem_resp_bits_xcpt_if;
  assign T336 = id_interrupt | io_imem_resp_bits_xcpt_ma;
  assign T337 = T338 & io_imem_resp_valid;
  assign T338 = id_interrupt & T339;
  assign T339 = take_pc_mem_wb ^ 1'h1;
  assign T340 = T342 & T341;
  assign T341 = mem_reg_replay_next ^ 1'h1;
  assign T342 = T343 & ex_reg_xcpt_interrupt;
  assign T343 = take_pc_mem_wb ^ 1'h1;
  assign killm_common = T347 | T344;
  assign T344 = mem_reg_valid ^ 1'h1;
  assign T345 = ctrl_killx ? 1'h0 : ex_reg_valid;
  assign T346 = ctrl_killd ? 1'h0 : 1'h1;
  assign T347 = T348 | mem_reg_xcpt;
  assign T348 = dcache_kill_mem | take_pc_wb;
  assign dcache_kill_mem = mem_reg_wen & io_dmem_replay_next_valid;
  assign T349 = ctrl_killx ? 1'h0 : ex_reg_wen;
  assign T350 = ctrl_killd ? 1'h0 : T351;
  assign T351 = T354 | T352;
  assign T352 = T353 == 32'h0;
  assign T353 = io_dpath_inst & 32'h28;
  assign T354 = T357 | T355;
  assign T355 = T356 == 32'h2010;
  assign T356 = io_dpath_inst & 32'h2010;
  assign T357 = T360 | T358;
  assign T358 = T359 == 32'h2008;
  assign T359 = io_dpath_inst & 32'h2008;
  assign T360 = T363 | T361;
  assign T361 = T362 == 32'h1010;
  assign T362 = io_dpath_inst & 32'h1010;
  assign T363 = T364 | T134;
  assign T364 = T367 | T365;
  assign T365 = T366 == 32'h10;
  assign T366 = io_dpath_inst & 32'h50;
  assign T367 = T368 == 32'h4;
  assign T368 = io_dpath_inst & 32'hc;
  assign T369 = wb_reg_div_mul_val | wb_dcache_miss;
  assign wb_dcache_miss = wb_reg_mem_val & T370;
  assign T370 = io_dmem_resp_valid ^ 1'h1;
  assign T371 = ctrl_killm ? 1'h0 : mem_reg_mem_val;
  assign T372 = ctrl_killm ? 1'h0 : mem_reg_div_mul_val;
  assign T373 = ex_reg_div_mul_val & io_dpath_div_mul_rdy;
  assign T374 = ctrl_killd ? 1'h0 : T375;
  assign T375 = T378 | T376;
  assign T376 = T377 == 32'h2004020;
  assign T377 = io_dpath_inst & 32'h2004064;
  assign T378 = T379 == 32'h2000030;
  assign T379 = io_dpath_inst & 32'h2004074;
  assign T380 = io_dpath_ll_wen | T125;
  assign id_wen_not0 = T351 & T381;
  assign T381 = T112 != 5'h0;
  assign T382 = T400 | T383;
  assign T383 = id_renx2_not0 & T384;
  assign T384 = T390 & T385;
  assign T385 = T386 - 1'h1;
  assign T386 = 1'h1 << T387;
  assign T387 = T388 + 5'h1;
  assign T388 = T389 - T389;
  assign T389 = io_dpath_inst[5'h18:5'h14];
  assign T390 = T114 >> T389;
  assign id_renx2_not0 = T392 & T391;
  assign T391 = T389 != 5'h0;
  assign T392 = T395 | T393;
  assign T393 = T394 == 32'h20;
  assign T394 = io_dpath_inst & 32'h34;
  assign T395 = T398 | T396;
  assign T396 = T397 == 32'h20;
  assign T397 = io_dpath_inst & 32'h64;
  assign T398 = T399 == 32'h20;
  assign T399 = io_dpath_inst & 32'h70;
  assign T400 = id_renx1_not0 & T401;
  assign T401 = T406 & T402;
  assign T402 = T403 - 1'h1;
  assign T403 = 1'h1 << T404;
  assign T404 = T405 + 5'h1;
  assign T405 = T29 - T29;
  assign T406 = T114 >> T29;
  assign id_renx1_not0 = T408 & T407;
  assign T407 = T29 != 5'h0;
  assign T408 = T411 | T409;
  assign T409 = T410 == 32'h2000;
  assign T410 = io_dpath_inst & 32'h2050;
  assign T411 = T414 | T412;
  assign T412 = T413 == 32'h2000;
  assign T413 = io_dpath_inst & 32'h6004;
  assign T414 = T417 | T415;
  assign T415 = T416 == 32'h1000;
  assign T416 = io_dpath_inst & 32'h5004;
  assign T417 = T420 | T418;
  assign T418 = T419 == 32'h0;
  assign T419 = io_dpath_inst & 32'h18;
  assign T420 = T421 == 32'h0;
  assign T421 = io_dpath_inst & 32'h44;
  assign T422 = T451 | id_wb_hazard;
  assign id_wb_hazard = T441 | T423;
  assign T423 = fp_data_hazard_wb & T424;
  assign T424 = wb_dcache_miss | wb_reg_fp_val;
  assign T425 = ctrl_killm ? 1'h0 : mem_reg_fp_val;
  assign fp_data_hazard_wb = wb_reg_fp_wen & T426;
  assign T426 = T429 | T427;
  assign T427 = io_fpu_dec_wen & T428;
  assign T428 = T112 == io_dpath_wb_waddr;
  assign T429 = T433 | T430;
  assign T430 = io_fpu_dec_ren3 & T431;
  assign T431 = T432 == io_dpath_wb_waddr;
  assign T432 = io_dpath_inst[5'h1f:5'h1b];
  assign T433 = T436 | T434;
  assign T434 = io_fpu_dec_ren2 & T435;
  assign T435 = T389 == io_dpath_wb_waddr;
  assign T436 = io_fpu_dec_ren1 & T437;
  assign T437 = T29 == io_dpath_wb_waddr;
  assign T438 = ctrl_killm ? 1'h0 : mem_reg_fp_wen;
  assign T439 = ctrl_killx ? 1'h0 : ex_reg_fp_wen;
  assign T440 = ctrl_killd ? 1'h0 : 1'h0;
  assign T441 = data_hazard_wb & wb_set_sboard;
  assign data_hazard_wb = wb_reg_wen & T442;
  assign T442 = T445 | T443;
  assign T443 = id_wen_not0 & T444;
  assign T444 = T112 == io_dpath_wb_waddr;
  assign T445 = T448 | T446;
  assign T446 = id_renx2_not0 & T447;
  assign T447 = T389 == io_dpath_wb_waddr;
  assign T448 = id_renx1_not0 & T449;
  assign T449 = T29 == io_dpath_wb_waddr;
  assign T450 = ctrl_killm ? 1'h0 : mem_reg_wen;
  assign T451 = id_ex_hazard | id_mem_hazard;
  assign id_mem_hazard = T464 | T452;
  assign T452 = fp_data_hazard_mem & mem_reg_fp_val;
  assign fp_data_hazard_mem = mem_reg_fp_wen & T453;
  assign T453 = T456 | T454;
  assign T454 = io_fpu_dec_wen & T455;
  assign T455 = T112 == io_dpath_mem_waddr;
  assign T456 = T459 | T457;
  assign T457 = io_fpu_dec_ren3 & T458;
  assign T458 = T432 == io_dpath_mem_waddr;
  assign T459 = T462 | T460;
  assign T460 = io_fpu_dec_ren2 & T461;
  assign T461 = T389 == io_dpath_mem_waddr;
  assign T462 = io_fpu_dec_ren1 & T463;
  assign T463 = T29 == io_dpath_mem_waddr;
  assign T464 = data_hazard_mem & T465;
  assign T465 = T466 | mem_reg_rocc_val;
  assign T466 = T467 | mem_reg_fp_val;
  assign T467 = T468 | mem_reg_div_mul_val;
  assign T468 = T517 | T469;
  assign T469 = mem_reg_mem_val & mem_reg_slow_bypass;
  assign T470 = T516 ? ex_slow_bypass : mem_reg_slow_bypass;
  assign ex_slow_bypass = T489 | T471;
  assign T471 = T484 | T472;
  assign T472 = 3'h5 == ex_reg_mem_type;
  assign T473 = T483 ? T474 : ex_reg_mem_type;
  assign T474 = T475;
  assign T475 = {T481, T476};
  assign T476 = {T479, T477};
  assign T477 = T478 == 32'h1000;
  assign T478 = io_dpath_inst & 32'h1000;
  assign T479 = T480 == 32'h2000;
  assign T480 = io_dpath_inst & 32'h2000;
  assign T481 = T482 == 32'h4000;
  assign T482 = io_dpath_inst & 32'h4000;
  assign T483 = ctrl_killd ^ 1'h1;
  assign T484 = T486 | T485;
  assign T485 = 3'h1 == ex_reg_mem_type;
  assign T486 = T488 | T487;
  assign T487 = 3'h4 == ex_reg_mem_type;
  assign T488 = 3'h0 == ex_reg_mem_type;
  assign T489 = ex_reg_mem_cmd == 5'h7;
  assign T490 = T483 ? T491 : ex_reg_mem_cmd;
  assign T491 = {1'h0, T492};
  assign T492 = {T514, T493};
  assign T493 = {T508, T494};
  assign T494 = {T503, T495};
  assign T495 = T498 | T496;
  assign T496 = T497 == 32'h20000020;
  assign T497 = io_dpath_inst & 32'h20000020;
  assign T498 = T501 | T499;
  assign T499 = T500 == 32'h18000020;
  assign T500 = io_dpath_inst & 32'h18000020;
  assign T501 = T502 == 32'h20;
  assign T502 = io_dpath_inst & 32'h28;
  assign T503 = T506 | T504;
  assign T504 = T505 == 32'h40000008;
  assign T505 = io_dpath_inst & 32'h40000008;
  assign T506 = T507 == 32'h10000008;
  assign T507 = io_dpath_inst & 32'h10000008;
  assign T508 = T511 | T509;
  assign T509 = T510 == 32'h80000008;
  assign T510 = io_dpath_inst & 32'h80000008;
  assign T511 = T512 | T506;
  assign T512 = T513 == 32'h8000008;
  assign T513 = io_dpath_inst & 32'h8000008;
  assign T514 = T515 == 32'h8;
  assign T515 = io_dpath_inst & 32'h18000008;
  assign T516 = ctrl_killx ^ 1'h1;
  assign T517 = mem_reg_csr != 2'h0;
  assign T518 = ctrl_killx ? 2'h0 : ex_reg_csr;
  assign T519 = ctrl_killd ? 2'h0 : T22;
  assign data_hazard_mem = mem_reg_wen & T520;
  assign T520 = T523 | T521;
  assign T521 = id_wen_not0 & T522;
  assign T522 = T112 == io_dpath_mem_waddr;
  assign T523 = T526 | T524;
  assign T524 = id_renx2_not0 & T525;
  assign T525 = T389 == io_dpath_mem_waddr;
  assign T526 = id_renx1_not0 & T527;
  assign T527 = T29 == io_dpath_mem_waddr;
  assign id_ex_hazard = T541 | T528;
  assign T528 = fp_data_hazard_ex & T529;
  assign T529 = ex_reg_mem_val | ex_reg_fp_val;
  assign fp_data_hazard_ex = ex_reg_fp_wen & T530;
  assign T530 = T533 | T531;
  assign T531 = io_fpu_dec_wen & T532;
  assign T532 = T112 == io_dpath_ex_waddr;
  assign T533 = T536 | T534;
  assign T534 = io_fpu_dec_ren3 & T535;
  assign T535 = T432 == io_dpath_ex_waddr;
  assign T536 = T539 | T537;
  assign T537 = io_fpu_dec_ren2 & T538;
  assign T538 = T389 == io_dpath_ex_waddr;
  assign T539 = io_fpu_dec_ren1 & T540;
  assign T540 = T29 == io_dpath_ex_waddr;
  assign T541 = data_hazard_ex & T542;
  assign T542 = T543 | ex_reg_rocc_val;
  assign T543 = T544 | ex_reg_fp_val;
  assign T544 = T545 | ex_reg_div_mul_val;
  assign T545 = T546 | ex_reg_mem_val;
  assign T546 = T547 | ex_reg_jalr;
  assign T547 = ex_reg_csr != 2'h0;
  assign data_hazard_ex = ex_reg_wen & T548;
  assign T548 = T551 | T549;
  assign T549 = id_wen_not0 & T550;
  assign T550 = T112 == io_dpath_ex_waddr;
  assign T551 = T554 | T552;
  assign T552 = id_renx2_not0 & T553;
  assign T553 = T389 == io_dpath_ex_waddr;
  assign T554 = id_renx1_not0 & T555;
  assign T555 = T29 == io_dpath_ex_waddr;
  assign T556 = T557 | take_pc_mem_wb;
  assign T557 = io_imem_resp_valid ^ 1'h1;
  assign T558 = wb_dcache_miss & ex_reg_load_use;
  assign T559 = ctrl_killd ? 1'h0 : id_load_use;
  assign id_load_use = T560;
  assign T560 = mem_reg_mem_val & T561;
  assign T561 = data_hazard_mem | fp_data_hazard_mem;
  assign replay_ex_structural = T564 | T562;
  assign T562 = ex_reg_div_mul_val & T563;
  assign T563 = io_dpath_div_mul_rdy ^ 1'h1;
  assign T564 = ex_reg_mem_val & T565;
  assign T565 = io_dmem_req_ready ^ 1'h1;
  assign T566 = take_pc_mem_wb ^ 1'h1;
  assign T567 = ctrl_killx ? 1'h0 : ex_reg_sret;
  assign T568 = ctrl_killd ? 1'h0 : T167;
  assign T569 = replay_wb | wb_reg_xcpt;
  assign replay_wb = replay_wb_common | T570;
  assign T570 = wb_reg_rocc_val & T571;
  assign T571 = io_rocc_cmd_ready ^ 1'h1;
  assign replay_wb_common = T572 | io_dpath_csr_replay;
  assign T572 = io_dmem_resp_bits_nack | wb_reg_replay;
  assign T573 = replay_mem & T574;
  assign T574 = take_pc_wb ^ 1'h1;
  assign replay_mem = T575 | fpu_kill_mem;
  assign T575 = dcache_kill_mem | mem_reg_replay;
  assign io_rocc_s = io_dpath_status_s;
  assign io_rocc_cmd_valid = wb_rocc_val;
  assign wb_rocc_val = wb_reg_rocc_val & T576;
  assign T576 = replay_wb_common ^ 1'h1;
  assign io_fpu_killm = killm_common;
  assign io_fpu_killx = ctrl_killx;
  assign io_fpu_valid = 1'h0;
  assign io_dmem_req_bits_cmd = ex_reg_mem_cmd;
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_req_bits_typ = ex_reg_mem_type;
  assign io_dmem_req_bits_kill = T577;
  assign T577 = killm_common | mem_xcpt;
  assign io_dmem_req_valid = ex_reg_mem_val;
  assign io_imem_invalidate = wb_reg_flush_inst;
  assign T578 = ctrl_killm ? 1'h0 : mem_reg_flush_inst;
  assign T579 = ctrl_killx ? 1'h0 : ex_reg_flush_inst;
  assign T580 = ctrl_killd ? 1'h0 : T98;
  assign io_imem_btb_update_bits_incorrectTarget = take_pc_mem;
  assign io_imem_btb_update_bits_isReturn = T581;
  assign T581 = mem_reg_jalr & io_dpath_mem_rs1_ra;
  assign io_imem_btb_update_bits_isCall = T582;
  assign T582 = mem_reg_wen & T583;
  assign T583 = io_dpath_mem_waddr[1'h0:1'h0];
  assign io_imem_btb_update_bits_isJump = T584;
  assign T584 = mem_reg_jal | mem_reg_jalr;
  assign io_imem_btb_update_bits_taken = T585;
  assign T585 = mem_reg_jal | T586;
  assign T586 = mem_reg_branch & io_dpath_mem_br_taken;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign T587 = T590 ? ex_reg_btb_resp_bht_value : mem_reg_btb_resp_bht_value;
  assign T588 = T589 ? io_imem_btb_resp_bits_bht_value : ex_reg_btb_resp_bht_value;
  assign T589 = T483 & io_imem_btb_resp_valid;
  assign T590 = T516 & ex_reg_btb_hit;
  assign T591 = ctrl_killd ? 1'h0 : io_imem_btb_resp_valid;
  assign io_imem_btb_update_bits_prediction_bits_bht_index = mem_reg_btb_resp_bht_index;
  assign T592 = T590 ? ex_reg_btb_resp_bht_index : mem_reg_btb_resp_bht_index;
  assign T593 = T589 ? io_imem_btb_resp_bits_bht_index : ex_reg_btb_resp_bht_index;
  assign io_imem_btb_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign T594 = T590 ? ex_reg_btb_resp_entry : mem_reg_btb_resp_entry;
  assign T595 = T589 ? io_imem_btb_resp_bits_entry : ex_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign T596 = T590 ? ex_reg_btb_resp_target : mem_reg_btb_resp_target;
  assign T597 = T589 ? io_imem_btb_resp_bits_target : ex_reg_btb_resp_target;
  assign io_imem_btb_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign T598 = T590 ? ex_reg_btb_resp_taken : mem_reg_btb_resp_taken;
  assign T599 = T589 ? io_imem_btb_resp_bits_taken : ex_reg_btb_resp_taken;
  assign io_imem_btb_update_bits_prediction_valid = mem_reg_btb_hit;
  assign T600 = T516 ? ex_reg_btb_hit : mem_reg_btb_hit;
  assign io_imem_btb_update_valid = T601;
  assign T601 = T602 | mem_reg_jalr;
  assign T602 = mem_reg_branch | mem_reg_jal;
  assign io_imem_resp_ready = T603;
  assign T603 = T604 | ctrl_draind;
  assign T604 = ctrl_stalld ^ 1'h1;
  assign io_imem_req_valid = take_pc_mem_wb;
  assign io_dpath_badvaddr_wen = wb_reg_xcpt;
  assign io_dpath_cause = wb_reg_cause;
  assign T605 = mem_xcpt ? mem_cause : wb_reg_cause;
  assign mem_cause = T157 ? mem_reg_cause : T606;
  assign T606 = {60'h0, T607};
  assign T607 = T156 ? 4'h8 : T608;
  assign T608 = T154 ? 4'h9 : T609;
  assign T609 = T152 ? 4'ha : 4'hb;
  assign T610 = ex_xcpt ? ex_cause : mem_reg_cause;
  assign ex_cause = T160 ? ex_reg_cause : 64'h2;
  assign T611 = id_xcpt ? id_cause : ex_reg_cause;
  assign id_cause = id_interrupt ? id_interrupt_cause : T612;
  assign T612 = {60'h0, T613};
  assign T613 = io_imem_resp_bits_xcpt_ma ? 4'h0 : T614;
  assign T614 = io_imem_resp_bits_xcpt_if ? 4'h1 : T615;
  assign T615 = T191 ? 4'h2 : T616;
  assign T616 = id_csr_privileged ? 4'h3 : T617;
  assign T617 = T165 ? 4'h3 : T618;
  assign T618 = T162 ? 4'h6 : 4'hc;
  assign id_interrupt_cause = T61 ? 64'h8000000000000000 : T619;
  assign T619 = T58 ? 64'h8000000000000001 : T620;
  assign T620 = T54 ? 64'h8000000000000002 : T621;
  assign T621 = T50 ? 64'h8000000000000003 : T622;
  assign T622 = T46 ? 64'h8000000000000004 : T623;
  assign T623 = T42 ? 64'h8000000000000005 : T624;
  assign T624 = T38 ? 64'h8000000000000006 : 64'h8000000000000007;
  assign io_dpath_exception = wb_reg_xcpt;
  assign io_dpath_retire = T625;
  assign T625 = wb_reg_valid & T626;
  assign T626 = replay_wb ^ 1'h1;
  assign T627 = ctrl_killm ? 1'h0 : mem_reg_valid;
  assign io_dpath_ll_ready = T628;
  assign T628 = wb_reg_wen ^ 1'h1;
  assign io_dpath_bypass_src_0 = T629;
  assign T629 = T638 ? 2'h0 : T630;
  assign T630 = T636 ? 2'h1 : T631;
  assign T631 = T632 ? 2'h2 : 2'h3;
  assign T632 = T634 & T633;
  assign T633 = io_dpath_mem_waddr == T29;
  assign T634 = mem_reg_wen & T635;
  assign T635 = mem_reg_mem_val ^ 1'h1;
  assign T636 = ex_reg_wen & T637;
  assign T637 = io_dpath_ex_waddr == T29;
  assign T638 = 5'h0 == T29;
  assign io_dpath_bypass_src_1 = T639;
  assign T639 = T646 ? 2'h0 : T640;
  assign T640 = T644 ? 2'h1 : T641;
  assign T641 = T642 ? 2'h2 : 2'h3;
  assign T642 = T634 & T643;
  assign T643 = io_dpath_mem_waddr == T389;
  assign T644 = ex_reg_wen & T645;
  assign T645 = io_dpath_ex_waddr == T389;
  assign T646 = 5'h0 == T389;
  assign io_dpath_bypass_0 = T647;
  assign T647 = T650 | T648;
  assign T648 = mem_reg_wen & T649;
  assign T649 = io_dpath_mem_waddr == T29;
  assign T650 = T651 | T632;
  assign T651 = T638 | T636;
  assign io_dpath_bypass_1 = T652;
  assign T652 = T655 | T653;
  assign T653 = mem_reg_wen & T654;
  assign T654 = io_dpath_mem_waddr == T389;
  assign T655 = T656 | T642;
  assign T656 = T646 | T644;
  assign io_dpath_mem_rocc_val = mem_reg_rocc_val;
  assign io_dpath_ex_rocc_val = ex_reg_rocc_val;
  assign io_dpath_ex_rs2_val = T657;
  assign T657 = T658 | ex_reg_rocc_val;
  assign T658 = ex_reg_mem_val & T659;
  assign T659 = T663 | T660;
  assign T660 = T662 | T661;
  assign T661 = ex_reg_mem_cmd == 5'h4;
  assign T662 = ex_reg_mem_cmd[2'h3:2'h3];
  assign T663 = T665 | T664;
  assign T664 = ex_reg_mem_cmd == 5'h7;
  assign T665 = ex_reg_mem_cmd == 5'h1;
  assign io_dpath_ex_mem_type = ex_reg_mem_type;
  assign io_dpath_wb_wen = T666;
  assign T666 = wb_reg_wen & T667;
  assign T667 = replay_wb ^ 1'h1;
  assign io_dpath_mem_wen = mem_reg_wen;
  assign io_dpath_mem_branch = mem_reg_branch;
  assign io_dpath_mem_jalr = mem_reg_jalr;
  assign io_dpath_ex_valid = ex_reg_valid;
  assign io_dpath_ex_wen = ex_reg_wen;
  assign io_dpath_mem_fp_val = mem_reg_fp_val;
  assign io_dpath_ex_fp_val = ex_reg_fp_val;
  assign io_dpath_wb_load = T668;
  assign T668 = wb_reg_mem_val & wb_reg_wen;
  assign io_dpath_mem_load = T669;
  assign T669 = mem_reg_mem_val & mem_reg_wen;
  assign io_dpath_sret = wb_reg_sret;
  assign io_dpath_csr = T670;
  assign T670 = {1'h0, wb_reg_csr};
  assign T671 = ctrl_killm ? 2'h0 : mem_reg_csr;
  assign io_dpath_div_mul_kill = T672;
  assign T672 = mem_reg_div_mul_val & killm_common;
  assign io_dpath_div_mul_val = ex_reg_div_mul_val;
  assign io_dpath_fn_alu = T673;
  assign T673 = T674;
  assign T674 = {T710, T675};
  assign T675 = {T699, T676};
  assign T676 = {T685, T677};
  assign T677 = T680 | T678;
  assign T678 = T679 == 32'h7000;
  assign T679 = io_dpath_inst & 32'h7044;
  assign T680 = T683 | T681;
  assign T681 = T682 == 32'h1040;
  assign T682 = io_dpath_inst & 32'h1058;
  assign T683 = T684 == 32'h1010;
  assign T684 = io_dpath_inst & 32'h3054;
  assign T685 = T688 | T686;
  assign T686 = T687 == 32'h40001010;
  assign T687 = io_dpath_inst & 32'h40001054;
  assign T688 = T691 | T689;
  assign T689 = T690 == 32'h40000030;
  assign T690 = io_dpath_inst & 32'h40003034;
  assign T691 = T694 | T692;
  assign T692 = T693 == 32'h6010;
  assign T693 = io_dpath_inst & 32'h6054;
  assign T694 = T697 | T695;
  assign T695 = T696 == 32'h3010;
  assign T696 = io_dpath_inst & 32'h3054;
  assign T697 = T698 == 32'h2040;
  assign T698 = io_dpath_inst & 32'h2058;
  assign T699 = T702 | T700;
  assign T700 = T701 == 32'h4040;
  assign T701 = io_dpath_inst & 32'h4058;
  assign T702 = T705 | T703;
  assign T703 = T704 == 32'h4010;
  assign T704 = io_dpath_inst & 32'h5054;
  assign T705 = T708 | T706;
  assign T706 = T707 == 32'h4010;
  assign T707 = io_dpath_inst & 32'h40004054;
  assign T708 = T709 == 32'h2010;
  assign T709 = io_dpath_inst & 32'h2054;
  assign T710 = T713 | T711;
  assign T711 = T712 == 32'h40001010;
  assign T712 = io_dpath_inst & 32'h40003054;
  assign T713 = T714 | T689;
  assign T714 = T143 | T715;
  assign T715 = T716 == 32'h2010;
  assign T716 = io_dpath_inst & 32'h6054;
  assign io_dpath_fn_dw = T717;
  assign T717 = T718;
  assign T718 = T721 | T719;
  assign T719 = T720 == 32'h0;
  assign T720 = io_dpath_inst & 32'h8;
  assign T721 = T722 == 32'h0;
  assign T722 = io_dpath_inst & 32'h10;
  assign io_dpath_sel_imm = T723;
  assign T723 = T724;
  assign T724 = {T734, T725};
  assign T725 = {T731, T726};
  assign T726 = T729 | T727;
  assign T727 = T728 == 32'h40;
  assign T728 = io_dpath_inst & 32'h44;
  assign T729 = T730 == 32'h8;
  assign T730 = io_dpath_inst & 32'h18;
  assign T731 = T732 | T729;
  assign T732 = T733 == 32'h4;
  assign T733 = io_dpath_inst & 32'h44;
  assign T734 = T737 | T735;
  assign T735 = T736 == 32'h10;
  assign T736 = io_dpath_inst & 32'h14;
  assign T737 = T738 | T139;
  assign T738 = T739 == 32'h0;
  assign T739 = io_dpath_inst & 32'h24;
  assign io_dpath_sel_alu1 = T740;
  assign T740 = T741;
  assign T741 = {T749, T742};
  assign T742 = T743 | T418;
  assign T743 = T744 | T420;
  assign T744 = T747 | T745;
  assign T745 = T746 == 32'h0;
  assign T746 = io_dpath_inst & 32'h50;
  assign T747 = T748 == 32'h0;
  assign T748 = io_dpath_inst & 32'h4004;
  assign T749 = T750 | T134;
  assign T750 = T751 == 32'h4;
  assign T751 = io_dpath_inst & 32'h24;
  assign io_dpath_sel_alu2 = T752;
  assign T752 = {1'h0, T753};
  assign T753 = T754;
  assign T754 = {T765, T755};
  assign T755 = T758 | T756;
  assign T756 = T757 == 32'h4050;
  assign T757 = io_dpath_inst & 32'h4050;
  assign T758 = T759 | T134;
  assign T759 = T760 | T367;
  assign T760 = T763 | T761;
  assign T761 = T762 == 32'h0;
  assign T762 = io_dpath_inst & 32'h20;
  assign T763 = T764 == 32'h0;
  assign T764 = io_dpath_inst & 32'h58;
  assign T765 = T768 | T766;
  assign T766 = T767 == 32'h4000;
  assign T767 = io_dpath_inst & 32'h4008;
  assign T768 = T769 | T418;
  assign T769 = T770 | T420;
  assign T770 = T771 == 32'h0;
  assign T771 = io_dpath_inst & 32'h48;
  assign io_dpath_ren_0 = T408;
  assign io_dpath_ren_1 = T392;
  assign io_dpath_killd = T772;
  assign T772 = take_pc_mem_wb | T773;
  assign T773 = ctrl_stalld & T774;
  assign T774 = ctrl_draind ^ 1'h1;
  assign io_dpath_sel_pc = T775;
  assign T775 = {1'h0, T776};
  assign T776 = wb_reg_xcpt ? 2'h3 : T777;
  assign T777 = wb_reg_sret ? 2'h3 : T778;
  assign T778 = replay_wb ? 2'h2 : 2'h1;

  always @(posedge clk) begin
    wb_reg_xcpt <= T1;
    if(ctrl_killm) begin
      wb_reg_sret <= 1'h0;
    end else begin
      wb_reg_sret <= T5;
    end
    mem_reg_replay <= T7;
    if(ctrl_killx) begin
      mem_reg_replay_next <= 1'h0;
    end else begin
      mem_reg_replay_next <= ex_reg_replay_next;
    end
    if(ctrl_killd) begin
      ex_reg_replay_next <= 1'h0;
    end else begin
      ex_reg_replay_next <= T10;
    end
    if(reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      id_reg_fence <= T86;
    end
    if(ctrl_killd) begin
      ex_reg_mem_val <= 1'h0;
    end else begin
      ex_reg_mem_val <= T89;
    end
    if(reset) begin
      R118 <= 32'h0;
    end else if(T380) begin
      R118 <= T122;
    end else if(io_dpath_ll_wen) begin
      R118 <= T114;
    end
    if(ctrl_killm) begin
      wb_reg_rocc_val <= 1'h0;
    end else begin
      wb_reg_rocc_val <= mem_reg_rocc_val;
    end
    if(ctrl_killx) begin
      mem_reg_rocc_val <= 1'h0;
    end else begin
      mem_reg_rocc_val <= ex_reg_rocc_val;
    end
    if(ctrl_killd) begin
      ex_reg_rocc_val <= 1'h0;
    end else begin
      ex_reg_rocc_val <= T129;
    end
    if(ctrl_killx) begin
      mem_reg_jal <= 1'h0;
    end else begin
      mem_reg_jal <= ex_reg_jal;
    end
    if(ctrl_killd) begin
      ex_reg_jal <= 1'h0;
    end else begin
      ex_reg_jal <= T134;
    end
    if(ctrl_killx) begin
      mem_reg_jalr <= 1'h0;
    end else begin
      mem_reg_jalr <= ex_reg_jalr;
    end
    if(ctrl_killd) begin
      ex_reg_jalr <= 1'h0;
    end else begin
      ex_reg_jalr <= T139;
    end
    if(ctrl_killx) begin
      mem_reg_branch <= 1'h0;
    end else begin
      mem_reg_branch <= ex_reg_branch;
    end
    if(ctrl_killd) begin
      ex_reg_branch <= 1'h0;
    end else begin
      ex_reg_branch <= T143;
    end
    if(ctrl_killx) begin
      mem_reg_fp_val <= 1'h0;
    end else begin
      mem_reg_fp_val <= ex_reg_fp_val;
    end
    if(ctrl_killd) begin
      ex_reg_fp_val <= 1'h0;
    end else begin
      ex_reg_fp_val <= 1'h0;
    end
    if(ctrl_killx) begin
      mem_reg_mem_val <= 1'h0;
    end else begin
      mem_reg_mem_val <= ex_reg_mem_val;
    end
    if(ctrl_killx) begin
      mem_reg_xcpt <= 1'h0;
    end else begin
      mem_reg_xcpt <= ex_xcpt;
    end
    if(ctrl_killd) begin
      ex_reg_xcpt <= 1'h0;
    end else begin
      ex_reg_xcpt <= id_xcpt;
    end
    ex_reg_xcpt_interrupt <= T337;
    mem_reg_xcpt_interrupt <= T340;
    if(ctrl_killx) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= ex_reg_valid;
    end
    if(ctrl_killd) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= 1'h1;
    end
    if(ctrl_killx) begin
      mem_reg_wen <= 1'h0;
    end else begin
      mem_reg_wen <= ex_reg_wen;
    end
    if(ctrl_killd) begin
      ex_reg_wen <= 1'h0;
    end else begin
      ex_reg_wen <= T351;
    end
    if(ctrl_killm) begin
      wb_reg_mem_val <= 1'h0;
    end else begin
      wb_reg_mem_val <= mem_reg_mem_val;
    end
    if(ctrl_killm) begin
      wb_reg_div_mul_val <= 1'h0;
    end else begin
      wb_reg_div_mul_val <= mem_reg_div_mul_val;
    end
    mem_reg_div_mul_val <= T373;
    if(ctrl_killd) begin
      ex_reg_div_mul_val <= 1'h0;
    end else begin
      ex_reg_div_mul_val <= T375;
    end
    if(ctrl_killm) begin
      wb_reg_fp_val <= 1'h0;
    end else begin
      wb_reg_fp_val <= mem_reg_fp_val;
    end
    if(ctrl_killm) begin
      wb_reg_fp_wen <= 1'h0;
    end else begin
      wb_reg_fp_wen <= mem_reg_fp_wen;
    end
    if(ctrl_killx) begin
      mem_reg_fp_wen <= 1'h0;
    end else begin
      mem_reg_fp_wen <= ex_reg_fp_wen;
    end
    if(ctrl_killd) begin
      ex_reg_fp_wen <= 1'h0;
    end else begin
      ex_reg_fp_wen <= 1'h0;
    end
    if(ctrl_killm) begin
      wb_reg_wen <= 1'h0;
    end else begin
      wb_reg_wen <= mem_reg_wen;
    end
    if(T516) begin
      mem_reg_slow_bypass <= ex_slow_bypass;
    end
    if(T483) begin
      ex_reg_mem_type <= T474;
    end
    if(T483) begin
      ex_reg_mem_cmd <= T491;
    end
    if(ctrl_killx) begin
      mem_reg_csr <= 2'h0;
    end else begin
      mem_reg_csr <= ex_reg_csr;
    end
    if(ctrl_killd) begin
      ex_reg_csr <= 2'h0;
    end else begin
      ex_reg_csr <= T22;
    end
    if(ctrl_killd) begin
      ex_reg_load_use <= 1'h0;
    end else begin
      ex_reg_load_use <= id_load_use;
    end
    if(ctrl_killx) begin
      mem_reg_sret <= 1'h0;
    end else begin
      mem_reg_sret <= ex_reg_sret;
    end
    if(ctrl_killd) begin
      ex_reg_sret <= 1'h0;
    end else begin
      ex_reg_sret <= T167;
    end
    wb_reg_replay <= T573;
    if(ctrl_killm) begin
      wb_reg_flush_inst <= 1'h0;
    end else begin
      wb_reg_flush_inst <= mem_reg_flush_inst;
    end
    if(ctrl_killx) begin
      mem_reg_flush_inst <= 1'h0;
    end else begin
      mem_reg_flush_inst <= ex_reg_flush_inst;
    end
    if(ctrl_killd) begin
      ex_reg_flush_inst <= 1'h0;
    end else begin
      ex_reg_flush_inst <= T98;
    end
    if(T590) begin
      mem_reg_btb_resp_bht_value <= ex_reg_btb_resp_bht_value;
    end
    if(T589) begin
      ex_reg_btb_resp_bht_value <= io_imem_btb_resp_bits_bht_value;
    end
    if(ctrl_killd) begin
      ex_reg_btb_hit <= 1'h0;
    end else begin
      ex_reg_btb_hit <= io_imem_btb_resp_valid;
    end
    if(T590) begin
      mem_reg_btb_resp_bht_index <= ex_reg_btb_resp_bht_index;
    end
    if(T589) begin
      ex_reg_btb_resp_bht_index <= io_imem_btb_resp_bits_bht_index;
    end
    if(T590) begin
      mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
    end
    if(T589) begin
      ex_reg_btb_resp_entry <= io_imem_btb_resp_bits_entry;
    end
    if(T590) begin
      mem_reg_btb_resp_target <= ex_reg_btb_resp_target;
    end
    if(T589) begin
      ex_reg_btb_resp_target <= io_imem_btb_resp_bits_target;
    end
    if(T590) begin
      mem_reg_btb_resp_taken <= ex_reg_btb_resp_taken;
    end
    if(T589) begin
      ex_reg_btb_resp_taken <= io_imem_btb_resp_bits_taken;
    end
    if(T516) begin
      mem_reg_btb_hit <= ex_reg_btb_hit;
    end
    if(mem_xcpt) begin
      wb_reg_cause <= mem_cause;
    end
    if(ex_xcpt) begin
      mem_reg_cause <= ex_cause;
    end
    if(id_xcpt) begin
      ex_reg_cause <= id_cause;
    end
    if(ctrl_killm) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= mem_reg_valid;
    end
    if(ctrl_killm) begin
      wb_reg_csr <= 2'h0;
    end else begin
      wb_reg_csr <= mem_reg_csr;
    end
  end
endmodule

module ALU(
    input  io_dw,
    input [3:0] io_fn,
    input [63:0] io_in2,
    input [63:0] io_in1,
    output[63:0] io_out,
    output[63:0] io_adder_out
);

  wire[63:0] sum;
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire[63:0] T3;
  wire[63:0] T4;
  wire[31:0] T5;
  wire[63:0] out64;
  wire[63:0] T6;
  wire[63:0] T7;
  wire[63:0] T8;
  wire[63:0] T9;
  wire[63:0] T10;
  wire[63:0] T11;
  wire cmp;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[63:0] T26;
  wire T27;
  wire[63:0] T28;
  wire T29;
  wire[63:0] T30;
  wire T31;
  wire[63:0] shout_l;
  wire[63:0] T32;
  wire[63:0] T33;
  wire[62:0] T34;
  wire[63:0] T35;
  wire[63:0] T36;
  wire[63:0] T37;
  wire[61:0] T38;
  wire[63:0] T39;
  wire[63:0] T40;
  wire[63:0] T41;
  wire[59:0] T42;
  wire[63:0] T43;
  wire[63:0] T44;
  wire[63:0] T45;
  wire[55:0] T46;
  wire[63:0] T47;
  wire[63:0] T48;
  wire[63:0] T49;
  wire[47:0] T50;
  wire[63:0] T51;
  wire[63:0] T52;
  wire[63:0] T53;
  wire[31:0] T54;
  wire[63:0] T55;
  wire[64:0] T56;
  wire[5:0] shamt;
  wire[5:0] T57;
  wire[4:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[64:0] T62;
  wire[64:0] T63;
  wire[63:0] shin;
  wire[63:0] T64;
  wire[63:0] T65;
  wire[63:0] T66;
  wire[62:0] T67;
  wire[63:0] T68;
  wire[63:0] T69;
  wire[63:0] T70;
  wire[61:0] T71;
  wire[63:0] T72;
  wire[63:0] T73;
  wire[63:0] T74;
  wire[59:0] T75;
  wire[63:0] T76;
  wire[63:0] T77;
  wire[63:0] T78;
  wire[55:0] T79;
  wire[63:0] T80;
  wire[63:0] T81;
  wire[63:0] T82;
  wire[47:0] T83;
  wire[63:0] T84;
  wire[63:0] T85;
  wire[63:0] T86;
  wire[31:0] T87;
  wire[63:0] shin_r;
  wire[31:0] T88;
  wire[31:0] shin_hi;
  wire[31:0] shin_hi_32;
  wire[31:0] T89;
  wire[31:0] T90;
  wire T91;
  wire T92;
  wire[31:0] T93;
  wire T94;
  wire[63:0] T95;
  wire[63:0] T96;
  wire[31:0] T97;
  wire[63:0] T98;
  wire[63:0] T99;
  wire[47:0] T100;
  wire[63:0] T101;
  wire[63:0] T102;
  wire[55:0] T103;
  wire[63:0] T104;
  wire[63:0] T105;
  wire[59:0] T106;
  wire[63:0] T107;
  wire[63:0] T108;
  wire[61:0] T109;
  wire[63:0] T110;
  wire[63:0] T111;
  wire[62:0] T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire[63:0] T119;
  wire[63:0] T120;
  wire[31:0] T121;
  wire[63:0] T122;
  wire[63:0] T123;
  wire[47:0] T124;
  wire[63:0] T125;
  wire[63:0] T126;
  wire[55:0] T127;
  wire[63:0] T128;
  wire[63:0] T129;
  wire[59:0] T130;
  wire[63:0] T131;
  wire[63:0] T132;
  wire[61:0] T133;
  wire[63:0] T134;
  wire[63:0] T135;
  wire[62:0] T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire[31:0] out_hi;
  wire[31:0] T144;
  wire[31:0] T145;
  wire T146;
  wire[31:0] T147;
  wire T148;


  assign io_adder_out = sum;
  assign sum = io_in1 + T0;
  assign T0 = T2 ? T1 : io_in2;
  assign T1 = 64'h0 - io_in2;
  assign T2 = io_fn[2'h3:2'h3];
  assign io_out = T3;
  assign T3 = T4;
  assign T4 = {out_hi, T5};
  assign T5 = out64[5'h1f:1'h0];
  assign out64 = T141 ? sum : T6;
  assign T6 = T138 ? T55 : T7;
  assign T7 = T137 ? shout_l : T8;
  assign T8 = T31 ? T30 : T9;
  assign T9 = T29 ? T28 : T10;
  assign T10 = T27 ? T26 : T11;
  assign T11 = {63'h0, cmp};
  assign cmp = T25 ^ T12;
  assign T12 = T23 ? T22 : T13;
  assign T13 = T19 ? T18 : T14;
  assign T14 = T17 ? T16 : T15;
  assign T15 = io_in1[6'h3f:6'h3f];
  assign T16 = io_in2[6'h3f:6'h3f];
  assign T17 = io_fn[1'h1:1'h1];
  assign T18 = sum[6'h3f:6'h3f];
  assign T19 = T21 == T20;
  assign T20 = io_in2[6'h3f:6'h3f];
  assign T21 = io_in1[6'h3f:6'h3f];
  assign T22 = sum == 64'h0;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_fn[2'h2:2'h2];
  assign T25 = io_fn[1'h0:1'h0];
  assign T26 = io_in1 ^ io_in2;
  assign T27 = io_fn == 4'h4;
  assign T28 = io_in1 | io_in2;
  assign T29 = io_fn == 4'h6;
  assign T30 = io_in1 & io_in2;
  assign T31 = io_fn == 4'h7;
  assign shout_l = T134 | T32;
  assign T32 = T33 & 64'haaaaaaaaaaaaaaaa;
  assign T33 = T34 << 1'h1;
  assign T34 = T35[6'h3e:1'h0];
  assign T35 = T131 | T36;
  assign T36 = T37 & 64'hcccccccccccccccc;
  assign T37 = T38 << 2'h2;
  assign T38 = T39[6'h3d:1'h0];
  assign T39 = T128 | T40;
  assign T40 = T41 & 64'hf0f0f0f0f0f0f0f0;
  assign T41 = T42 << 3'h4;
  assign T42 = T43[6'h3b:1'h0];
  assign T43 = T125 | T44;
  assign T44 = T45 & 64'hff00ff00ff00ff00;
  assign T45 = T46 << 4'h8;
  assign T46 = T47[6'h37:1'h0];
  assign T47 = T122 | T48;
  assign T48 = T49 & 64'hffff0000ffff0000;
  assign T49 = T50 << 5'h10;
  assign T50 = T51[6'h2f:1'h0];
  assign T51 = T119 | T52;
  assign T52 = T53 & 64'hffffffff00000000;
  assign T53 = T54 << 6'h20;
  assign T54 = T55[5'h1f:1'h0];
  assign T55 = T56[6'h3f:1'h0];
  assign T56 = $signed(T62) >>> shamt;
  assign shamt = T57;
  assign T57 = {T59, T58};
  assign T58 = io_in2[3'h4:1'h0];
  assign T59 = T61 & T60;
  assign T60 = io_dw == 1'h1;
  assign T61 = io_in2[3'h5:3'h5];
  assign T62 = T63;
  assign T63 = {T116, shin};
  assign shin = T113 ? shin_r : T64;
  assign T64 = T110 | T65;
  assign T65 = T66 & 64'haaaaaaaaaaaaaaaa;
  assign T66 = T67 << 1'h1;
  assign T67 = T68[6'h3e:1'h0];
  assign T68 = T107 | T69;
  assign T69 = T70 & 64'hcccccccccccccccc;
  assign T70 = T71 << 2'h2;
  assign T71 = T72[6'h3d:1'h0];
  assign T72 = T104 | T73;
  assign T73 = T74 & 64'hf0f0f0f0f0f0f0f0;
  assign T74 = T75 << 3'h4;
  assign T75 = T76[6'h3b:1'h0];
  assign T76 = T101 | T77;
  assign T77 = T78 & 64'hff00ff00ff00ff00;
  assign T78 = T79 << 4'h8;
  assign T79 = T80[6'h37:1'h0];
  assign T80 = T98 | T81;
  assign T81 = T82 & 64'hffff0000ffff0000;
  assign T82 = T83 << 5'h10;
  assign T83 = T84[6'h2f:1'h0];
  assign T84 = T95 | T85;
  assign T85 = T86 & 64'hffffffff00000000;
  assign T86 = T87 << 6'h20;
  assign T87 = shin_r[5'h1f:1'h0];
  assign shin_r = {shin_hi, T88};
  assign T88 = io_in1[5'h1f:1'h0];
  assign shin_hi = T94 ? T93 : shin_hi_32;
  assign shin_hi_32 = T92 ? T89 : 32'h0;
  assign T89 = 32'h0 - T90;
  assign T90 = {31'h0, T91};
  assign T91 = io_in1[5'h1f:5'h1f];
  assign T92 = io_fn[2'h3:2'h3];
  assign T93 = io_in1[6'h3f:6'h20];
  assign T94 = io_dw == 1'h1;
  assign T95 = T96 & 64'hffffffff;
  assign T96 = {32'h0, T97};
  assign T97 = shin_r >> 6'h20;
  assign T98 = T99 & 64'hffff0000ffff;
  assign T99 = {16'h0, T100};
  assign T100 = T84 >> 5'h10;
  assign T101 = T102 & 64'hff00ff00ff00ff;
  assign T102 = {8'h0, T103};
  assign T103 = T80 >> 4'h8;
  assign T104 = T105 & 64'hf0f0f0f0f0f0f0f;
  assign T105 = {4'h0, T106};
  assign T106 = T76 >> 3'h4;
  assign T107 = T108 & 64'h3333333333333333;
  assign T108 = {2'h0, T109};
  assign T109 = T72 >> 2'h2;
  assign T110 = T111 & 64'h5555555555555555;
  assign T111 = {1'h0, T112};
  assign T112 = T68 >> 1'h1;
  assign T113 = T115 | T114;
  assign T114 = io_fn == 4'hb;
  assign T115 = io_fn == 4'h5;
  assign T116 = T118 & T117;
  assign T117 = shin[6'h3f:6'h3f];
  assign T118 = io_fn[2'h3:2'h3];
  assign T119 = T120 & 64'hffffffff;
  assign T120 = {32'h0, T121};
  assign T121 = T55 >> 6'h20;
  assign T122 = T123 & 64'hffff0000ffff;
  assign T123 = {16'h0, T124};
  assign T124 = T51 >> 5'h10;
  assign T125 = T126 & 64'hff00ff00ff00ff;
  assign T126 = {8'h0, T127};
  assign T127 = T47 >> 4'h8;
  assign T128 = T129 & 64'hf0f0f0f0f0f0f0f;
  assign T129 = {4'h0, T130};
  assign T130 = T43 >> 3'h4;
  assign T131 = T132 & 64'h3333333333333333;
  assign T132 = {2'h0, T133};
  assign T133 = T39 >> 2'h2;
  assign T134 = T135 & 64'h5555555555555555;
  assign T135 = {1'h0, T136};
  assign T136 = T35 >> 1'h1;
  assign T137 = io_fn == 4'h1;
  assign T138 = T140 | T139;
  assign T139 = io_fn == 4'hb;
  assign T140 = io_fn == 4'h5;
  assign T141 = T143 | T142;
  assign T142 = io_fn == 4'ha;
  assign T143 = io_fn == 4'h0;
  assign out_hi = T148 ? T147 : T144;
  assign T144 = 32'h0 - T145;
  assign T145 = {31'h0, T146};
  assign T146 = out64[5'h1f:5'h1f];
  assign T147 = out64[6'h3f:6'h20];
  assign T148 = io_dw == 1'h1;
endmodule

module MulDiv(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [3:0] io_req_bits_fn,
    input  io_req_bits_dw,
    input [63:0] io_req_bits_in1,
    input [63:0] io_req_bits_in2,
    input [4:0] io_req_bits_tag,
    input  io_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[63:0] io_resp_bits_data,
    output[4:0] io_resp_bits_tag
);

  reg [4:0] req_tag;
  wire[4:0] T0;
  wire T1;
  wire[63:0] T2;
  wire[63:0] T3;
  reg [129:0] remainder;
  wire[129:0] T4;
  wire[129:0] T5;
  wire[129:0] T6;
  wire[129:0] T7;
  wire[129:0] T8;
  wire[129:0] T9;
  wire[129:0] T10;
  wire[63:0] negated_remainder;
  wire[63:0] T11;
  wire T12;
  wire T13;
  reg  isMul;
  wire T14;
  wire T15;
  wire T16;
  wire[3:0] T17;
  wire T18;
  wire[3:0] T19;
  wire T20;
  wire T21;
  reg [2:0] state;
  wire[2:0] T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire T30;
  wire[2:0] T31;
  reg  neg_out;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  reg  isHi;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire[3:0] T41;
  wire T42;
  wire[3:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire[64:0] subtractor;
  reg [64:0] divisor;
  wire[64:0] T47;
  wire[64:0] T48;
  wire T49;
  wire T50;
  wire T51;
  wire[64:0] T52;
  wire[63:0] rhs_in;
  wire[31:0] T53;
  wire[31:0] T54;
  wire[31:0] T55;
  wire[31:0] T56;
  wire rhs_sign;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[3:0] T63;
  wire[31:0] T64;
  wire T65;
  wire[64:0] T66;
  wire T67;
  reg [6:0] count;
  wire[6:0] T68;
  wire[6:0] T69;
  wire[6:0] T70;
  wire[6:0] T71;
  wire T72;
  wire T73;
  wire[6:0] T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire lhs_sign;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire[3:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire[2:0] T91;
  wire T92;
  wire T93;
  wire[2:0] T94;
  wire[2:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire[2:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire[129:0] T104;
  wire[129:0] T105;
  wire[63:0] T106;
  wire[129:0] T107;
  wire[129:0] T108;
  wire[64:0] T109;
  wire[63:0] T110;
  wire[128:0] T111;
  wire[63:0] T112;
  wire[128:0] T113;
  wire[128:0] T114;
  wire[62:0] T115;
  wire[63:0] T116;
  wire[128:0] T117;
  wire[63:0] T118;
  wire[64:0] T119;
  wire[65:0] T120;
  wire[65:0] T121;
  wire[64:0] T122;
  wire[64:0] T123;
  wire T124;
  wire[65:0] T125;
  wire[1:0] T126;
  wire[1:0] T127;
  wire T128;
  wire[64:0] T129;
  wire[64:0] T130;
  wire[64:0] T131;
  wire[129:0] T132;
  wire[128:0] T133;
  wire[64:0] T134;
  wire T135;
  wire[63:0] T136;
  wire[63:0] T137;
  wire[63:0] T138;
  wire[63:0] T139;
  wire[129:0] T140;
  wire[63:0] lhs_in;
  wire[31:0] T141;
  wire[31:0] T142;
  wire[31:0] T143;
  wire[31:0] T144;
  wire[31:0] T145;
  wire T146;
  wire[63:0] T147;
  wire[31:0] T148;
  wire[31:0] T149;
  wire[31:0] T150;
  wire T151;
  wire T152;
  reg  req_dw;
  wire T153;
  wire T154;
  wire T155;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    req_tag = {1{$random}};
    remainder = {5{$random}};
    isMul = {1{$random}};
    state = {1{$random}};
    neg_out = {1{$random}};
    isHi = {1{$random}};
    divisor = {3{$random}};
    count = {1{$random}};
    req_dw = {1{$random}};
  end
`endif

  assign io_resp_bits_tag = req_tag;
  assign T0 = T1 ? io_req_bits_tag : req_tag;
  assign T1 = io_req_ready & io_req_valid;
  assign io_resp_bits_data = T2;
  assign T2 = T152 ? T147 : T3;
  assign T3 = remainder[6'h3f:1'h0];
  assign T4 = T1 ? T140 : T5;
  assign T5 = T75 ? T132 : T6;
  assign T6 = T72 ? T107 : T7;
  assign T7 = T90 ? T105 : T8;
  assign T8 = T30 ? T104 : T9;
  assign T9 = T12 ? T10 : remainder;
  assign T10 = {66'h0, negated_remainder};
  assign negated_remainder = 64'h0 - T11;
  assign T11 = remainder[6'h3f:1'h0];
  assign T12 = T21 & T13;
  assign T13 = T20 | isMul;
  assign T14 = T1 ? T15 : isMul;
  assign T15 = T18 | T16;
  assign T16 = T17 == 4'h8;
  assign T17 = io_req_bits_fn & 4'h8;
  assign T18 = T19 == 4'h0;
  assign T19 = io_req_bits_fn & 4'h4;
  assign T20 = remainder[6'h3f:6'h3f];
  assign T21 = state == 3'h1;
  assign T22 = reset ? 3'h0 : T23;
  assign T23 = T1 ? T100 : T24;
  assign T24 = T98 ? 3'h0 : T25;
  assign T25 = T96 ? T94 : T26;
  assign T26 = T92 ? T91 : T27;
  assign T27 = T90 ? T31 : T28;
  assign T28 = T30 ? 3'h5 : T29;
  assign T29 = T21 ? 3'h2 : state;
  assign T30 = state == 3'h4;
  assign T31 = neg_out ? 3'h4 : 3'h5;
  assign T32 = T1 ? T78 : T33;
  assign T33 = T34 ? 1'h0 : neg_out;
  assign T34 = T75 & T35;
  assign T35 = T44 & T36;
  assign T36 = isHi ^ 1'h1;
  assign T37 = T1 ? T38 : isHi;
  assign T38 = T39 | T16;
  assign T39 = T42 | T40;
  assign T40 = T41 == 4'h2;
  assign T41 = io_req_bits_fn & 4'h2;
  assign T42 = T43 == 4'h1;
  assign T43 = io_req_bits_fn & 4'h5;
  assign T44 = T67 & T45;
  assign T45 = T46 ^ 1'h1;
  assign T46 = subtractor[7'h40:7'h40];
  assign subtractor = T66 - divisor;
  assign T47 = T1 ? T52 : T48;
  assign T48 = T49 ? subtractor : divisor;
  assign T49 = T21 & T50;
  assign T50 = T51 | isMul;
  assign T51 = divisor[6'h3f:6'h3f];
  assign T52 = {rhs_sign, rhs_in};
  assign rhs_in = {T54, T53};
  assign T53 = io_req_bits_in2[5'h1f:1'h0];
  assign T54 = T65 ? T64 : T55;
  assign T55 = 32'h0 - T56;
  assign T56 = {31'h0, rhs_sign};
  assign rhs_sign = T61 & T57;
  assign T57 = T60 ? T59 : T58;
  assign T58 = io_req_bits_in2[5'h1f:5'h1f];
  assign T59 = io_req_bits_in2[6'h3f:6'h3f];
  assign T60 = io_req_bits_dw == 1'h1;
  assign T61 = T62 | T18;
  assign T62 = T63 == 4'h0;
  assign T63 = io_req_bits_fn & 4'h9;
  assign T64 = io_req_bits_in2[6'h3f:6'h20];
  assign T65 = io_req_bits_dw == 1'h1;
  assign T66 = remainder[8'h80:7'h40];
  assign T67 = count == 7'h0;
  assign T68 = T1 ? 7'h0 : T69;
  assign T69 = T75 ? T74 : T70;
  assign T70 = T72 ? T71 : count;
  assign T71 = count + 7'h1;
  assign T72 = T73 & isMul;
  assign T73 = state == 3'h2;
  assign T74 = count + 7'h1;
  assign T75 = T77 & T76;
  assign T76 = isMul ^ 1'h1;
  assign T77 = state == 3'h2;
  assign T78 = T89 & T79;
  assign T79 = T38 ? lhs_sign : T80;
  assign T80 = lhs_sign != rhs_sign;
  assign lhs_sign = T85 & T81;
  assign T81 = T84 ? T83 : T82;
  assign T82 = io_req_bits_in1[5'h1f:5'h1f];
  assign T83 = io_req_bits_in1[6'h3f:6'h3f];
  assign T84 = io_req_bits_dw == 1'h1;
  assign T85 = T88 | T86;
  assign T86 = T87 == 4'h0;
  assign T87 = io_req_bits_fn & 4'h3;
  assign T88 = T62 | T18;
  assign T89 = T15 ^ 1'h1;
  assign T90 = state == 3'h3;
  assign T91 = isHi ? 3'h3 : 3'h5;
  assign T92 = T72 & T93;
  assign T93 = count == 7'h3f;
  assign T94 = isHi ? 3'h3 : T95;
  assign T95 = neg_out ? 3'h4 : 3'h5;
  assign T96 = T75 & T97;
  assign T97 = count == 7'h40;
  assign T98 = T99 | io_kill;
  assign T99 = io_resp_ready & io_resp_valid;
  assign T100 = T101 ? 3'h1 : 3'h2;
  assign T101 = lhs_sign | T102;
  assign T102 = rhs_sign & T103;
  assign T103 = T15 ^ 1'h1;
  assign T104 = {66'h0, negated_remainder};
  assign T105 = {66'h0, T106};
  assign T106 = remainder[8'h80:7'h41];
  assign T107 = T108;
  assign T108 = {T131, T109};
  assign T109 = {1'h0, T110};
  assign T110 = T111[6'h3f:1'h0];
  assign T111 = {T130, T112};
  assign T112 = T113[6'h3f:1'h0];
  assign T113 = T114;
  assign T114 = {T120, T115};
  assign T115 = T116[6'h3f:1'h1];
  assign T116 = T117[6'h3f:1'h0];
  assign T117 = {T119, T118};
  assign T118 = remainder[6'h3f:1'h0];
  assign T119 = remainder[8'h81:7'h41];
  assign T120 = T125 + T121;
  assign T121 = {T124, T122};
  assign T122 = T123;
  assign T123 = T117[8'h80:7'h40];
  assign T124 = T122[7'h40:7'h40];
  assign T125 = $signed(T129) * $signed(T126);
  assign T126 = T127;
  assign T127 = {1'h0, T128};
  assign T128 = T116[1'h0:1'h0];
  assign T129 = divisor;
  assign T130 = T113[8'h80:7'h40];
  assign T131 = T111 >> 7'h40;
  assign T132 = {1'h0, T133};
  assign T133 = {T137, T134};
  assign T134 = {T136, T135};
  assign T135 = T46 ^ 1'h1;
  assign T136 = remainder[6'h3f:1'h0];
  assign T137 = T46 ? T139 : T138;
  assign T138 = subtractor[6'h3f:1'h0];
  assign T139 = remainder[7'h7f:7'h40];
  assign T140 = {66'h0, lhs_in};
  assign lhs_in = {T142, T141};
  assign T141 = io_req_bits_in1[5'h1f:1'h0];
  assign T142 = T146 ? T145 : T143;
  assign T143 = 32'h0 - T144;
  assign T144 = {31'h0, lhs_sign};
  assign T145 = io_req_bits_in1[6'h3f:6'h20];
  assign T146 = io_req_bits_dw == 1'h1;
  assign T147 = {T149, T148};
  assign T148 = remainder[5'h1f:1'h0];
  assign T149 = 32'h0 - T150;
  assign T150 = {31'h0, T151};
  assign T151 = remainder[5'h1f:5'h1f];
  assign T152 = req_dw == 1'h0;
  assign T153 = T1 ? io_req_bits_dw : req_dw;
  assign io_resp_valid = T154;
  assign T154 = state == 3'h5;
  assign io_req_ready = T155;
  assign T155 = state == 3'h0;

  always @(posedge clk) begin
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(T1) begin
      remainder <= T140;
    end else if(T75) begin
      remainder <= T132;
    end else if(T72) begin
      remainder <= T107;
    end else if(T90) begin
      remainder <= T105;
    end else if(T30) begin
      remainder <= T104;
    end else if(T12) begin
      remainder <= T10;
    end
    if(T1) begin
      isMul <= T15;
    end
    if(reset) begin
      state <= 3'h0;
    end else if(T1) begin
      state <= T100;
    end else if(T98) begin
      state <= 3'h0;
    end else if(T96) begin
      state <= T94;
    end else if(T92) begin
      state <= T91;
    end else if(T90) begin
      state <= T31;
    end else if(T30) begin
      state <= 3'h5;
    end else if(T21) begin
      state <= 3'h2;
    end
    if(T1) begin
      neg_out <= T78;
    end else if(T34) begin
      neg_out <= 1'h0;
    end
    if(T1) begin
      isHi <= T38;
    end
    if(T1) begin
      divisor <= T52;
    end else if(T49) begin
      divisor <= subtractor;
    end
    if(T1) begin
      count <= 7'h0;
    end else if(T75) begin
      count <= T74;
    end else if(T72) begin
      count <= T71;
    end
    if(T1) begin
      req_dw <= io_req_bits_dw;
    end
  end
endmodule

module CSRFile(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    input [11:0] io_rw_addr,
    input [1:0] io_rw_cmd,
    output[63:0] io_rw_rdata,
    input [63:0] io_rw_wdata,
    output[7:0] io_status_ip,
    output[7:0] io_status_im,
    output[6:0] io_status_zero,
    output io_status_er,
    output io_status_vm,
    output io_status_s64,
    output io_status_u64,
    output io_status_ef,
    output io_status_pei,
    output io_status_ei,
    output io_status_ps,
    output io_status_s,
    output[31:0] io_ptbr,
    output[43:0] io_evec,
    input  io_exception,
    input  io_retire,
    input [63:0] io_cause,
    input  io_badvaddr_wen,
    input [43:0] io_pc,
    input  io_sret,
    output io_fatc,
    output io_replay,
    output[63:0] io_time,
    output[2:0] io_fcsr_rm,
    input  io_fcsr_flags_valid,
    input [4:0] io_fcsr_flags_bits,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[3:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [3:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    //output io_rocc_exception
);

  reg [2:0] reg_frm;
  wire[2:0] T0;
  wire[63:0] T1;
  wire[63:0] T2;
  wire[63:0] T3;
  wire[63:0] wdata;
  reg [63:0] host_pcr_bits_data;
  wire[63:0] T4;
  wire[63:0] T5;
  wire T6;
  wire host_pcr_req_fire;
  wire T7;
  wire T8;
  reg  host_pcr_req_valid;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire[41:0] T13;
  wire[40:0] T14;
  wire[39:0] T15;
  wire[38:0] T16;
  wire[37:0] T17;
  wire[36:0] T18;
  wire[35:0] T19;
  wire[34:0] T20;
  wire[33:0] T21;
  wire[32:0] T22;
  wire[31:0] T23;
  wire[30:0] T24;
  wire[29:0] T25;
  wire[28:0] T26;
  wire[27:0] T27;
  wire[26:0] T28;
  wire[25:0] T29;
  wire[24:0] T30;
  wire[23:0] T31;
  wire[22:0] T32;
  wire[21:0] T33;
  wire[20:0] T34;
  wire[19:0] T35;
  wire[18:0] T36;
  wire[17:0] T37;
  wire[16:0] T38;
  wire[15:0] T39;
  wire[14:0] T40;
  wire[13:0] T41;
  wire[12:0] T42;
  wire[11:0] T43;
  wire[10:0] T44;
  wire[9:0] T45;
  wire[8:0] T46;
  wire[7:0] T47;
  wire[6:0] T48;
  wire[5:0] T49;
  wire[4:0] T50;
  wire[3:0] T51;
  wire[2:0] T52;
  wire[1:0] T53;
  wire T54;
  wire[11:0] T55;
  wire[11:0] addr;
  wire[11:0] T56;
  wire[10:0] T57;
  wire[10:0] T58;
  reg [4:0] host_pcr_bits_addr;
  wire[4:0] T59;
  wire T60;
  wire[11:0] T61;
  wire T62;
  wire[11:0] T63;
  wire T64;
  wire[11:0] T65;
  wire T66;
  wire[11:0] T67;
  wire T68;
  wire[11:0] T69;
  wire T70;
  wire[11:0] T71;
  wire T72;
  wire[11:0] T73;
  wire T74;
  wire[11:0] T75;
  wire T76;
  wire[11:0] T77;
  wire T78;
  wire[11:0] T79;
  wire T80;
  wire[11:0] T81;
  wire T82;
  wire[11:0] T83;
  wire T84;
  wire[11:0] T85;
  wire T86;
  wire[11:0] T87;
  wire T88;
  wire[11:0] T89;
  wire T90;
  wire[11:0] T91;
  wire T92;
  wire[11:0] T93;
  wire T94;
  wire[11:0] T95;
  wire T96;
  wire[11:0] T97;
  wire T98;
  wire[11:0] T99;
  wire T100;
  wire[11:0] T101;
  wire T102;
  wire[11:0] T103;
  wire T104;
  wire[11:0] T105;
  wire T106;
  wire[11:0] T107;
  wire T108;
  wire[11:0] T109;
  wire T110;
  wire[11:0] T111;
  wire T112;
  wire[11:0] T113;
  wire T114;
  wire[11:0] T115;
  wire T116;
  wire[11:0] T117;
  wire T118;
  wire[11:0] T119;
  wire T120;
  wire[11:0] T121;
  wire T122;
  wire[11:0] T123;
  wire T124;
  wire[11:0] T125;
  wire T126;
  wire[11:0] T127;
  wire T128;
  wire[11:0] T129;
  wire T130;
  wire[11:0] T131;
  wire T132;
  wire[11:0] T133;
  wire T134;
  wire[11:0] T135;
  wire T136;
  wire[11:0] T137;
  wire T138;
  wire[11:0] T139;
  wire T140;
  wire[11:0] T141;
  wire wen;
  wire T142;
  reg  host_pcr_bits_rw;
  wire T143;
  wire[63:0] T144;
  wire[58:0] T145;
  wire T146;
  wire T147;
  wire[63:0] T148;
  reg [5:0] R149;
  wire[5:0] T150;
  wire[5:0] T151;
  wire[5:0] T152;
  wire[6:0] T153;
  wire[6:0] T154;
  wire[5:0] T155;
  wire[63:0] T156;
  wire T157;
  wire T158;
  reg [57:0] R159;
  wire[57:0] T160;
  wire[57:0] T161;
  wire[57:0] T162;
  wire[57:0] T163;
  wire T164;
  wire[57:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire[43:0] T170;
  wire[43:0] T171;
  reg [43:0] reg_epc;
  wire[43:0] T172;
  wire[43:0] T173;
  wire[43:0] T174;
  wire[43:0] T175;
  wire[43:0] T176;
  wire T177;
  wire T178;
  wire[43:0] T179;
  wire[42:0] T180;
  reg [42:0] reg_evec;
  wire[42:0] T181;
  wire[42:0] T182;
  wire[42:0] T183;
  wire T184;
  wire T185;
  wire T186;
  reg [31:0] reg_ptbr;
  wire[31:0] T187;
  wire[31:0] T188;
  wire[31:0] T189;
  wire[18:0] T190;
  wire T191;
  wire T192;
  reg  reg_status_s;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  reg  reg_status_ps;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  reg  reg_status_ei;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  reg  reg_status_pei;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  reg  reg_status_ef;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  reg  reg_status_u64;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  reg  reg_status_s64;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  reg  reg_status_vm;
  wire T225;
  wire T226;
  wire T227;
  reg  reg_status_er;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  reg [6:0] reg_status_zero;
  wire[6:0] T232;
  wire[6:0] T233;
  wire[6:0] T234;
  wire[6:0] T235;
  reg [7:0] reg_status_im;
  wire[7:0] T236;
  wire[7:0] T237;
  wire[7:0] T238;
  wire[7:0] T239;
  wire[3:0] T240;
  wire[1:0] T241;
  reg  r_irq_ipi;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[1:0] T248;
  wire T249;
  reg [63:0] reg_fromhost;
  wire[63:0] T250;
  wire[63:0] T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  reg  r_irq_timer;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  reg [31:0] reg_compare;
  wire[31:0] T262;
  wire[31:0] T263;
  wire[31:0] T264;
  wire T265;
  wire T266;
  wire[31:0] T267;
  wire[63:0] T268;
  wire[63:0] T269;
  wire[63:0] T270;
  wire[63:0] T271;
  reg [63:0] reg_tohost;
  wire[63:0] T272;
  wire[63:0] T273;
  wire[63:0] T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire[63:0] T283;
  wire[63:0] T284;
  wire T285;
  reg  reg_stats;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire[63:0] T291;
  wire[63:0] T292;
  wire[1:0] T293;
  wire[63:0] T294;
  wire[63:0] T295;
  wire[1:0] T296;
  wire T297;
  wire[63:0] T298;
  wire[63:0] T299;
  wire[1:0] T300;
  wire[63:0] T301;
  wire[63:0] T302;
  wire[1:0] T303;
  wire T304;
  wire[63:0] T305;
  wire[63:0] T306;
  wire T307;
  wire T308;
  wire[63:0] T309;
  wire[63:0] T310;
  wire[31:0] T311;
  wire[31:0] T312;
  wire[31:0] T313;
  wire[5:0] T314;
  wire[2:0] T315;
  wire[1:0] T316;
  wire[2:0] T317;
  wire[1:0] T318;
  wire[25:0] T319;
  wire[2:0] T320;
  wire[1:0] T321;
  wire[22:0] T322;
  wire[14:0] T323;
  wire[63:0] T324;
  wire[63:0] T325;
  reg [63:0] reg_cause;
  wire[63:0] T326;
  wire T327;
  wire[63:0] T328;
  wire[63:0] T329;
  wire[42:0] T330;
  wire[63:0] T331;
  wire[63:0] T332;
  wire[31:0] T333;
  wire[63:0] T334;
  wire[63:0] T335;
  wire[63:0] T336;
  wire[63:0] T337;
  wire[63:0] T338;
  wire[31:0] T339;
  wire[31:0] read_ptbr;
  wire[18:0] T340;
  wire[63:0] T341;
  wire[63:0] T342;
  wire[42:0] T343;
  reg [42:0] reg_badvaddr;
  wire[42:0] T344;
  wire[43:0] T345;
  wire[43:0] T346;
  wire[43:0] T347;
  wire[43:0] T348;
  wire[42:0] T349;
  wire T350;
  wire T351;
  wire[20:0] T352;
  wire T353;
  wire T354;
  wire[42:0] T355;
  wire T356;
  wire[63:0] T357;
  wire[63:0] T358;
  wire[43:0] T359;
  wire[63:0] T360;
  wire[63:0] T361;
  reg [63:0] reg_sup1;
  wire[63:0] T362;
  wire T363;
  wire T364;
  wire[63:0] T365;
  wire[63:0] T366;
  reg [63:0] reg_sup0;
  wire[63:0] T367;
  wire T368;
  wire T369;
  wire[63:0] T370;
  wire[63:0] T371;
  wire[63:0] T372;
  reg [5:0] R373;
  wire[5:0] T374;
  wire[5:0] T375;
  wire[5:0] T376;
  wire[6:0] T377;
  wire[6:0] T378;
  wire T379;
  reg [57:0] R380;
  wire[57:0] T381;
  wire[57:0] T382;
  wire[57:0] T383;
  wire T384;
  wire T385;
  wire T386;
  wire[63:0] T387;
  wire[63:0] T388;
  wire T389;
  wire[63:0] T390;
  wire[63:0] T391;
  wire T392;
  wire T393;
  wire T394;
  reg  host_pcr_rep_valid;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    reg_frm = {1{$random}};
    host_pcr_bits_data = {2{$random}};
    host_pcr_req_valid = {1{$random}};
    host_pcr_bits_addr = {1{$random}};
    host_pcr_bits_rw = {1{$random}};
    R149 = {1{$random}};
    R159 = {2{$random}};
    reg_epc = {2{$random}};
    reg_evec = {2{$random}};
    reg_ptbr = {1{$random}};
    reg_status_s = {1{$random}};
    reg_status_ps = {1{$random}};
    reg_status_ei = {1{$random}};
    reg_status_pei = {1{$random}};
    reg_status_ef = {1{$random}};
    reg_status_u64 = {1{$random}};
    reg_status_s64 = {1{$random}};
    reg_status_vm = {1{$random}};
    reg_status_er = {1{$random}};
    reg_status_zero = {1{$random}};
    reg_status_im = {1{$random}};
    r_irq_ipi = {1{$random}};
    reg_fromhost = {2{$random}};
    r_irq_timer = {1{$random}};
    reg_compare = {1{$random}};
    reg_tohost = {2{$random}};
    reg_stats = {1{$random}};
    reg_cause = {2{$random}};
    reg_badvaddr = {2{$random}};
    reg_sup1 = {2{$random}};
    reg_sup0 = {2{$random}};
    R373 = {1{$random}};
    R380 = {2{$random}};
    host_pcr_rep_valid = {1{$random}};
  end
`endif

  assign io_fcsr_rm = reg_frm;
  assign T0 = T1[2'h2:1'h0];
  assign T1 = T146 ? T144 : T2;
  assign T2 = T11 ? wdata : T3;
  assign T3 = {61'h0, reg_frm};
  assign wdata = T8 ? io_rw_wdata : host_pcr_bits_data;
  assign T4 = host_pcr_req_fire ? io_rw_rdata : T5;
  assign T5 = T6 ? io_host_pcr_req_bits_data : host_pcr_bits_data;
  assign T6 = io_host_pcr_req_ready & io_host_pcr_req_valid;
  assign host_pcr_req_fire = host_pcr_req_valid & T7;
  assign T7 = T8 ^ 1'h1;
  assign T8 = io_rw_cmd != 2'h0;
  assign T9 = host_pcr_req_fire ? 1'h0 : T10;
  assign T10 = T6 ? 1'h1 : host_pcr_req_valid;
  assign T11 = wen & T12;
  assign T12 = T13[1'h1:1'h1];
  assign T13 = {T140, T14};
  assign T14 = {T138, T15};
  assign T15 = {T136, T16};
  assign T16 = {T134, T17};
  assign T17 = {T132, T18};
  assign T18 = {T130, T19};
  assign T19 = {T128, T20};
  assign T20 = {T126, T21};
  assign T21 = {T124, T22};
  assign T22 = {T122, T23};
  assign T23 = {T120, T24};
  assign T24 = {T118, T25};
  assign T25 = {T116, T26};
  assign T26 = {T114, T27};
  assign T27 = {T112, T28};
  assign T28 = {T110, T29};
  assign T29 = {T108, T30};
  assign T30 = {T106, T31};
  assign T31 = {T104, T32};
  assign T32 = {T102, T33};
  assign T33 = {T100, T34};
  assign T34 = {T98, T35};
  assign T35 = {T96, T36};
  assign T36 = {T94, T37};
  assign T37 = {T92, T38};
  assign T38 = {T90, T39};
  assign T39 = {T88, T40};
  assign T40 = {T86, T41};
  assign T41 = {T84, T42};
  assign T42 = {T82, T43};
  assign T43 = {T80, T44};
  assign T44 = {T78, T45};
  assign T45 = {T76, T46};
  assign T46 = {T74, T47};
  assign T47 = {T72, T48};
  assign T48 = {T70, T49};
  assign T49 = {T68, T50};
  assign T50 = {T66, T51};
  assign T51 = {T64, T52};
  assign T52 = {T62, T53};
  assign T53 = {T60, T54};
  assign T54 = T55 == 12'h0;
  assign T55 = addr & 12'h482;
  assign addr = T8 ? io_rw_addr : T56;
  assign T56 = {1'h0, T57};
  assign T57 = T58 | 11'h500;
  assign T58 = {6'h0, host_pcr_bits_addr};
  assign T59 = T6 ? io_host_pcr_req_bits_addr : host_pcr_bits_addr;
  assign T60 = T61 == 12'h0;
  assign T61 = addr & 12'h481;
  assign T62 = T63 == 12'h3;
  assign T63 = addr & 12'h403;
  assign T64 = T65 == 12'h0;
  assign T65 = addr & 12'h403;
  assign T66 = T67 == 12'h0;
  assign T67 = addr & 12'h88f;
  assign T68 = T69 == 12'h401;
  assign T69 = addr & 12'hc0f;
  assign T70 = T71 == 12'h402;
  assign T71 = addr & 12'hc0f;
  assign T72 = T73 == 12'h403;
  assign T73 = addr & 12'hc0f;
  assign T74 = T75 == 12'h4;
  assign T75 = addr & 12'h80f;
  assign T76 = T77 == 12'h5;
  assign T77 = addr & 12'h80f;
  assign T78 = T79 == 12'h6;
  assign T79 = addr & 12'h80f;
  assign T80 = T81 == 12'h7;
  assign T81 = addr & 12'h80f;
  assign T82 = T83 == 12'h8;
  assign T83 = addr & 12'h80f;
  assign T84 = T85 == 12'h9;
  assign T85 = addr & 12'h80f;
  assign T86 = T87 == 12'ha;
  assign T87 = addr & 12'h80f;
  assign T88 = T89 == 12'hb;
  assign T89 = addr & 12'h80f;
  assign T90 = T91 == 12'hc;
  assign T91 = addr & 12'h80f;
  assign T92 = T93 == 12'hd;
  assign T93 = addr & 12'h81f;
  assign T94 = T95 == 12'he;
  assign T95 = addr & 12'h81f;
  assign T96 = T97 == 12'hf;
  assign T97 = addr & 12'h81f;
  assign T98 = T99 == 12'h10;
  assign T99 = addr & 12'h12;
  assign T100 = T101 == 12'h10;
  assign T101 = addr & 12'h11;
  assign T102 = T103 == 12'h13;
  assign T103 = addr & 12'h13;
  assign T104 = T105 == 12'h0;
  assign T105 = addr & 12'h183;
  assign T106 = T107 == 12'h801;
  assign T107 = addr & 12'h881;
  assign T108 = T109 == 12'h802;
  assign T109 = addr & 12'h882;
  assign T110 = T111 == 12'h880;
  assign T111 = addr & 12'h88f;
  assign T112 = T113 == 12'h81;
  assign T113 = addr & 12'h8f;
  assign T114 = T115 == 12'h82;
  assign T115 = addr & 12'h8f;
  assign T116 = T117 == 12'h803;
  assign T117 = addr & 12'h80f;
  assign T118 = T119 == 12'h4;
  assign T119 = addr & 12'h10f;
  assign T120 = T121 == 12'h5;
  assign T121 = addr & 12'h10f;
  assign T122 = T123 == 12'h6;
  assign T123 = addr & 12'h10f;
  assign T124 = T125 == 12'h7;
  assign T125 = addr & 12'h10f;
  assign T126 = T127 == 12'h8;
  assign T127 = addr & 12'h10f;
  assign T128 = T129 == 12'h9;
  assign T129 = addr & 12'h10f;
  assign T130 = T131 == 12'ha;
  assign T131 = addr & 12'h10f;
  assign T132 = T133 == 12'hb;
  assign T133 = addr & 12'h10f;
  assign T134 = T135 == 12'hc;
  assign T135 = addr & 12'h10f;
  assign T136 = T137 == 12'hd;
  assign T137 = addr & 12'h10f;
  assign T138 = T139 == 12'he;
  assign T139 = addr & 12'h10f;
  assign T140 = T141 == 12'hf;
  assign T141 = addr & 12'h10f;
  assign wen = T8 | T142;
  assign T142 = host_pcr_req_fire & host_pcr_bits_rw;
  assign T143 = T6 ? io_host_pcr_req_bits_rw : host_pcr_bits_rw;
  assign T144 = {5'h0, T145};
  assign T145 = wdata >> 3'h5;
  assign T146 = wen & T147;
  assign T147 = T13[2'h2:2'h2];
  assign io_time = T148;
  assign T148 = {R159, R149};
  assign T150 = reset ? 6'h0 : T151;
  assign T151 = T157 ? T155 : T152;
  assign T152 = T153[3'h5:1'h0];
  assign T153 = T154 + 7'h1;
  assign T154 = {1'h0, R149};
  assign T155 = T156[3'h5:1'h0];
  assign T156 = wdata;
  assign T157 = wen & T158;
  assign T158 = T13[4'ha:4'ha];
  assign T160 = reset ? 58'h0 : T161;
  assign T161 = T157 ? T165 : T162;
  assign T162 = T164 ? T163 : R159;
  assign T163 = R159 + 58'h1;
  assign T164 = T153[3'h6:3'h6];
  assign T165 = T156[6'h3f:3'h6];
  assign io_replay = T166;
  assign T166 = io_host_ipi_req_valid & T167;
  assign T167 = io_host_ipi_req_ready ^ 1'h1;
  assign io_fatc = T168;
  assign T168 = wen & T169;
  assign T169 = T13[5'h11:5'h11];
  assign io_evec = T170;
  assign T170 = T171;
  assign T171 = io_exception ? T179 : reg_epc;
  assign T172 = T177 ? T175 : T173;
  assign T173 = io_exception ? T174 : reg_epc;
  assign T174 = io_pc;
  assign T175 = T176;
  assign T176 = wdata[6'h2b:1'h0];
  assign T177 = wen & T178;
  assign T178 = T13[3'h6:3'h6];
  assign T179 = {T186, T180};
  assign T180 = reg_evec;
  assign T181 = T184 ? T182 : reg_evec;
  assign T182 = T183;
  assign T183 = wdata[6'h2a:1'h0];
  assign T184 = wen & T185;
  assign T185 = T13[4'hc:4'hc];
  assign T186 = T180[6'h2a:6'h2a];
  assign io_ptbr = reg_ptbr;
  assign T187 = T191 ? T188 : reg_ptbr;
  assign T188 = T189;
  assign T189 = {T190, 13'h0};
  assign T190 = wdata[5'h1f:4'hd];
  assign T191 = wen & T192;
  assign T192 = T13[4'h8:4'h8];
  assign io_status_s = reg_status_s;
  assign T193 = reset ? 1'h1 : T194;
  assign T194 = T201 ? T203 : T195;
  assign T195 = io_sret ? reg_status_ps : T196;
  assign T196 = io_exception ? 1'h1 : reg_status_s;
  assign T197 = reset ? 1'h0 : T198;
  assign T198 = T201 ? T200 : T199;
  assign T199 = io_exception ? reg_status_s : reg_status_ps;
  assign T200 = wdata[1'h1:1'h1];
  assign T201 = wen & T202;
  assign T202 = T13[4'he:4'he];
  assign T203 = wdata[1'h0:1'h0];
  assign io_status_ps = reg_status_ps;
  assign io_status_ei = reg_status_ei;
  assign T204 = reset ? 1'h0 : T205;
  assign T205 = T201 ? T212 : T206;
  assign T206 = io_sret ? reg_status_pei : T207;
  assign T207 = io_exception ? 1'h0 : reg_status_ei;
  assign T208 = reset ? 1'h0 : T209;
  assign T209 = T201 ? T211 : T210;
  assign T210 = io_exception ? reg_status_ei : reg_status_pei;
  assign T211 = wdata[2'h3:2'h3];
  assign T212 = wdata[2'h2:2'h2];
  assign io_status_pei = reg_status_pei;
  assign io_status_ef = reg_status_ef;
  assign T213 = reset ? 1'h0 : T214;
  assign T214 = T201 ? 1'h0 : T215;
  assign T215 = T201 ? T216 : reg_status_ef;
  assign T216 = wdata[3'h4:3'h4];
  assign io_status_u64 = reg_status_u64;
  assign T217 = reset ? 1'h1 : T218;
  assign T218 = T201 ? 1'h1 : T219;
  assign T219 = T201 ? T220 : reg_status_u64;
  assign T220 = wdata[3'h5:3'h5];
  assign io_status_s64 = reg_status_s64;
  assign T221 = reset ? 1'h1 : T222;
  assign T222 = T201 ? 1'h1 : T223;
  assign T223 = T201 ? T224 : reg_status_s64;
  assign T224 = wdata[3'h6:3'h6];
  assign io_status_vm = reg_status_vm;
  assign T225 = reset ? 1'h0 : T226;
  assign T226 = T201 ? T227 : reg_status_vm;
  assign T227 = wdata[3'h7:3'h7];
  assign io_status_er = reg_status_er;
  assign T228 = reset ? 1'h0 : T229;
  assign T229 = T201 ? 1'h0 : T230;
  assign T230 = T201 ? T231 : reg_status_er;
  assign T231 = wdata[4'h8:4'h8];
  assign io_status_zero = reg_status_zero;
  assign T232 = reset ? 7'h0 : T233;
  assign T233 = T201 ? 7'h0 : T234;
  assign T234 = T201 ? T235 : reg_status_zero;
  assign T235 = wdata[4'hf:4'h9];
  assign io_status_im = reg_status_im;
  assign T236 = reset ? 8'h0 : T237;
  assign T237 = T201 ? T238 : reg_status_im;
  assign T238 = wdata[5'h17:5'h10];
  assign io_status_ip = T239;
  assign T239 = {T240, 4'h0};
  assign T240 = {T248, T241};
  assign T241 = {r_irq_ipi, 1'h0};
  assign T242 = reset ? 1'h1 : T243;
  assign T243 = io_host_ipi_rep_valid ? 1'h1 : T244;
  assign T244 = T246 ? T245 : r_irq_ipi;
  assign T245 = wdata[1'h0:1'h0];
  assign T246 = wen & T247;
  assign T247 = T13[5'h13:5'h13];
  assign T248 = {r_irq_timer, T249};
  assign T249 = reg_fromhost != 64'h0;
  assign T250 = reset ? 64'h0 : T251;
  assign T251 = T252 ? wdata : reg_fromhost;
  assign T252 = T256 & T253;
  assign T253 = T255 | T254;
  assign T254 = host_pcr_req_fire ^ 1'h1;
  assign T255 = reg_fromhost == 64'h0;
  assign T256 = wen & T257;
  assign T257 = T13[5'h16:5'h16];
  assign T258 = reset ? 1'h0 : T259;
  assign T259 = T265 ? 1'h0 : T260;
  assign T260 = T261 ? 1'h1 : r_irq_timer;
  assign T261 = T267 == reg_compare;
  assign T262 = T265 ? T263 : reg_compare;
  assign T263 = T264;
  assign T264 = wdata[5'h1f:1'h0];
  assign T265 = wen & T266;
  assign T266 = T13[4'hb:4'hb];
  assign T267 = T148[5'h1f:1'h0];
  assign io_rw_rdata = T268;
  assign T268 = T270 | T269;
  assign T269 = T257 ? reg_fromhost : 64'h0;
  assign T270 = T283 | T271;
  assign T271 = T276 ? reg_tohost : 64'h0;
  assign T272 = reset ? 64'h0 : T273;
  assign T273 = T279 ? wdata : T274;
  assign T274 = T275 ? 64'h0 : reg_tohost;
  assign T275 = T277 & T276;
  assign T276 = T13[5'h15:5'h15];
  assign T277 = host_pcr_req_fire & T278;
  assign T278 = host_pcr_bits_rw ^ 1'h1;
  assign T279 = T282 & T280;
  assign T280 = T281 | host_pcr_req_fire;
  assign T281 = reg_tohost == 64'h0;
  assign T282 = wen & T276;
  assign T283 = T291 | T284;
  assign T284 = {63'h0, T285};
  assign T285 = T290 ? reg_stats : 1'h0;
  assign T286 = reset ? 1'h0 : T287;
  assign T287 = T289 ? T288 : reg_stats;
  assign T288 = wdata[1'h0:1'h0];
  assign T289 = wen & T290;
  assign T290 = T13[2'h3:2'h3];
  assign T291 = T294 | T292;
  assign T292 = {62'h0, T293};
  assign T293 = T247 ? 2'h2 : 2'h0;
  assign T294 = T298 | T295;
  assign T295 = {62'h0, T296};
  assign T296 = T297 ? 2'h2 : 2'h0;
  assign T297 = T13[5'h12:5'h12];
  assign T298 = T301 | T299;
  assign T299 = {62'h0, T300};
  assign T300 = T169 ? 2'h2 : 2'h0;
  assign T301 = T305 | T302;
  assign T302 = {62'h0, T303};
  assign T303 = T304 ? 2'h2 : 2'h0;
  assign T304 = T13[5'h10:5'h10];
  assign T305 = T309 | T306;
  assign T306 = {63'h0, T307};
  assign T307 = T308 ? io_host_id : 1'h0;
  assign T308 = T13[4'hf:4'hf];
  assign T309 = T324 | T310;
  assign T310 = {32'h0, T311};
  assign T311 = T202 ? T312 : 32'h0;
  assign T312 = T313;
  assign T313 = {T319, T314};
  assign T314 = {T317, T315};
  assign T315 = {io_status_ei, T316};
  assign T316 = {io_status_ps, io_status_s};
  assign T317 = {io_status_u64, T318};
  assign T318 = {io_status_ef, io_status_pei};
  assign T319 = {T322, T320};
  assign T320 = {io_status_er, T321};
  assign T321 = {io_status_vm, io_status_s64};
  assign T322 = {io_status_ip, T323};
  assign T323 = {io_status_im, io_status_zero};
  assign T324 = T328 | T325;
  assign T325 = T327 ? reg_cause : 64'h0;
  assign T326 = io_exception ? io_cause : reg_cause;
  assign T327 = T13[4'hd:4'hd];
  assign T328 = T331 | T329;
  assign T329 = {21'h0, T330};
  assign T330 = T185 ? reg_evec : 43'h0;
  assign T331 = T334 | T332;
  assign T332 = {32'h0, T333};
  assign T333 = T266 ? reg_compare : 32'h0;
  assign T334 = T336 | T335;
  assign T335 = T158 ? T148 : 64'h0;
  assign T336 = T337 | 64'h0;
  assign T337 = T341 | T338;
  assign T338 = {32'h0, T339};
  assign T339 = T192 ? read_ptbr : 32'h0;
  assign read_ptbr = T340 << 4'hd;
  assign T340 = reg_ptbr[5'h1f:4'hd];
  assign T341 = T357 | T342;
  assign T342 = {21'h0, T343};
  assign T343 = T356 ? reg_badvaddr : 43'h0;
  assign T344 = T345[6'h2a:1'h0];
  assign T345 = io_badvaddr_wen ? T347 : T346;
  assign T346 = {1'h0, reg_badvaddr};
  assign T347 = T348;
  assign T348 = {T350, T349};
  assign T349 = io_rw_wdata[6'h2a:1'h0];
  assign T350 = T354 ? T353 : T351;
  assign T351 = T352 != 21'h0;
  assign T352 = io_rw_wdata[6'h3f:6'h2b];
  assign T353 = T352 == 21'h1fffff;
  assign T354 = $signed(T355) < $signed(1'h0);
  assign T355 = T349;
  assign T356 = T13[3'h7:3'h7];
  assign T357 = T360 | T358;
  assign T358 = {20'h0, T359};
  assign T359 = T178 ? reg_epc : 44'h0;
  assign T360 = T365 | T361;
  assign T361 = T364 ? reg_sup1 : 64'h0;
  assign T362 = T363 ? wdata : reg_sup1;
  assign T363 = wen & T364;
  assign T364 = T13[3'h5:3'h5];
  assign T365 = T370 | T366;
  assign T366 = T369 ? reg_sup0 : 64'h0;
  assign T367 = T368 ? wdata : reg_sup0;
  assign T368 = wen & T369;
  assign T369 = T13[3'h4:3'h4];
  assign T370 = T387 | T371;
  assign T371 = T386 ? T372 : 64'h0;
  assign T372 = {R380, R373};
  assign T374 = reset ? 6'h0 : T375;
  assign T375 = T379 ? T376 : R373;
  assign T376 = T377[3'h5:1'h0];
  assign T377 = T378 + 7'h1;
  assign T378 = {1'h0, R373};
  assign T379 = io_retire != 1'h0;
  assign T381 = reset ? 58'h0 : T382;
  assign T382 = T384 ? T383 : R380;
  assign T383 = R380 + 58'h1;
  assign T384 = T379 & T385;
  assign T385 = T377[3'h6:3'h6];
  assign T386 = T13[5'h19:5'h19];
  assign T387 = T390 | T388;
  assign T388 = T389 ? T148 : 64'h0;
  assign T389 = T13[5'h18:5'h18];
  assign T390 = 64'h0 | T391;
  assign T391 = T392 ? T148 : 64'h0;
  assign T392 = T13[5'h17:5'h17];
  assign io_host_debug_stats_pcr = reg_stats;
  assign io_host_ipi_rep_ready = 1'h1;
  assign io_host_ipi_req_bits = T393;
  assign T393 = io_rw_wdata[1'h0:1'h0];
  assign io_host_ipi_req_valid = T394;
  assign T394 = T8 & T297;
  assign io_host_pcr_rep_bits = host_pcr_bits_data;
  assign io_host_pcr_rep_valid = host_pcr_rep_valid;
  assign T395 = T397 ? 1'h0 : T396;
  assign T396 = host_pcr_req_fire ? 1'h1 : host_pcr_rep_valid;
  assign T397 = io_host_pcr_rep_ready & io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = T398;
  assign T398 = T400 & T399;
  assign T399 = host_pcr_rep_valid ^ 1'h1;
  assign T400 = host_pcr_req_valid ^ 1'h1;

  always @(posedge clk) begin
    reg_frm <= T0;
    if(host_pcr_req_fire) begin
      host_pcr_bits_data <= io_rw_rdata;
    end else if(T6) begin
      host_pcr_bits_data <= io_host_pcr_req_bits_data;
    end
    if(host_pcr_req_fire) begin
      host_pcr_req_valid <= 1'h0;
    end else if(T6) begin
      host_pcr_req_valid <= 1'h1;
    end
    if(T6) begin
      host_pcr_bits_addr <= io_host_pcr_req_bits_addr;
    end
    if(T6) begin
      host_pcr_bits_rw <= io_host_pcr_req_bits_rw;
    end
    if(reset) begin
      R149 <= 6'h0;
    end else if(T157) begin
      R149 <= T155;
    end else begin
      R149 <= T152;
    end
    if(reset) begin
      R159 <= 58'h0;
    end else if(T157) begin
      R159 <= T165;
    end else if(T164) begin
      R159 <= T163;
    end
    if(T177) begin
      reg_epc <= T175;
    end else if(io_exception) begin
      reg_epc <= T174;
    end
    if(T184) begin
      reg_evec <= T182;
    end
    if(T191) begin
      reg_ptbr <= T188;
    end
    if(reset) begin
      reg_status_s <= 1'h1;
    end else if(T201) begin
      reg_status_s <= T203;
    end else if(io_sret) begin
      reg_status_s <= reg_status_ps;
    end else if(io_exception) begin
      reg_status_s <= 1'h1;
    end
    if(reset) begin
      reg_status_ps <= 1'h0;
    end else if(T201) begin
      reg_status_ps <= T200;
    end else if(io_exception) begin
      reg_status_ps <= reg_status_s;
    end
    if(reset) begin
      reg_status_ei <= 1'h0;
    end else if(T201) begin
      reg_status_ei <= T212;
    end else if(io_sret) begin
      reg_status_ei <= reg_status_pei;
    end else if(io_exception) begin
      reg_status_ei <= 1'h0;
    end
    if(reset) begin
      reg_status_pei <= 1'h0;
    end else if(T201) begin
      reg_status_pei <= T211;
    end else if(io_exception) begin
      reg_status_pei <= reg_status_ei;
    end
    if(reset) begin
      reg_status_ef <= 1'h0;
    end else if(T201) begin
      reg_status_ef <= 1'h0;
    end else if(T201) begin
      reg_status_ef <= T216;
    end
    if(reset) begin
      reg_status_u64 <= 1'h1;
    end else if(T201) begin
      reg_status_u64 <= 1'h1;
    end else if(T201) begin
      reg_status_u64 <= T220;
    end
    if(reset) begin
      reg_status_s64 <= 1'h1;
    end else if(T201) begin
      reg_status_s64 <= 1'h1;
    end else if(T201) begin
      reg_status_s64 <= T224;
    end
    if(reset) begin
      reg_status_vm <= 1'h0;
    end else if(T201) begin
      reg_status_vm <= T227;
    end
    if(reset) begin
      reg_status_er <= 1'h0;
    end else if(T201) begin
      reg_status_er <= 1'h0;
    end else if(T201) begin
      reg_status_er <= T231;
    end
    if(reset) begin
      reg_status_zero <= 7'h0;
    end else if(T201) begin
      reg_status_zero <= 7'h0;
    end else if(T201) begin
      reg_status_zero <= T235;
    end
    if(reset) begin
      reg_status_im <= 8'h0;
    end else if(T201) begin
      reg_status_im <= T238;
    end
    if(reset) begin
      r_irq_ipi <= 1'h1;
    end else if(io_host_ipi_rep_valid) begin
      r_irq_ipi <= 1'h1;
    end else if(T246) begin
      r_irq_ipi <= T245;
    end
    if(reset) begin
      reg_fromhost <= 64'h0;
    end else if(T252) begin
      reg_fromhost <= wdata;
    end
    if(reset) begin
      r_irq_timer <= 1'h0;
    end else if(T265) begin
      r_irq_timer <= 1'h0;
    end else if(T261) begin
      r_irq_timer <= 1'h1;
    end
    if(T265) begin
      reg_compare <= T263;
    end
    if(reset) begin
      reg_tohost <= 64'h0;
    end else if(T279) begin
      reg_tohost <= wdata;
    end else if(T275) begin
      reg_tohost <= 64'h0;
    end
    if(reset) begin
      reg_stats <= 1'h0;
    end else if(T289) begin
      reg_stats <= T288;
    end
    if(io_exception) begin
      reg_cause <= io_cause;
    end
    reg_badvaddr <= T344;
    if(T363) begin
      reg_sup1 <= wdata;
    end
    if(T368) begin
      reg_sup0 <= wdata;
    end
    if(reset) begin
      R373 <= 6'h0;
    end else if(T379) begin
      R373 <= T376;
    end
    if(reset) begin
      R380 <= 58'h0;
    end else if(T384) begin
      R380 <= T383;
    end
    if(T397) begin
      host_pcr_rep_valid <= 1'h0;
    end else if(host_pcr_req_fire) begin
      host_pcr_rep_valid <= 1'h1;
    end
  end
endmodule

module Datapath(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    input [2:0] io_ctrl_sel_pc,
    input  io_ctrl_killd,
    input  io_ctrl_ren_1,
    input  io_ctrl_ren_0,
    input [2:0] io_ctrl_sel_alu2,
    input [1:0] io_ctrl_sel_alu1,
    input [2:0] io_ctrl_sel_imm,
    input  io_ctrl_fn_dw,
    input [3:0] io_ctrl_fn_alu,
    input  io_ctrl_div_mul_val,
    input  io_ctrl_div_mul_kill,
    //input  io_ctrl_div_val
    //input  io_ctrl_div_kill
    input [2:0] io_ctrl_csr,
    input  io_ctrl_sret,
    input  io_ctrl_mem_load,
    input  io_ctrl_wb_load,
    input  io_ctrl_ex_fp_val,
    input  io_ctrl_mem_fp_val,
    input  io_ctrl_ex_wen,
    input  io_ctrl_ex_valid,
    input  io_ctrl_mem_jalr,
    input  io_ctrl_mem_branch,
    input  io_ctrl_mem_wen,
    input  io_ctrl_wb_wen,
    input [2:0] io_ctrl_ex_mem_type,
    input  io_ctrl_ex_rs2_val,
    input  io_ctrl_ex_rocc_val,
    input  io_ctrl_mem_rocc_val,
    input  io_ctrl_bypass_1,
    input  io_ctrl_bypass_0,
    input [1:0] io_ctrl_bypass_src_1,
    input [1:0] io_ctrl_bypass_src_0,
    input  io_ctrl_ll_ready,
    input  io_ctrl_retire,
    input  io_ctrl_exception,
    input [63:0] io_ctrl_cause,
    input  io_ctrl_badvaddr_wen,
    output[31:0] io_ctrl_inst,
    //output io_ctrl_jalr_eq
    output io_ctrl_mem_br_taken,
    output io_ctrl_mem_misprediction,
    output io_ctrl_div_mul_rdy,
    output io_ctrl_ll_wen,
    output[4:0] io_ctrl_ll_waddr,
    output[4:0] io_ctrl_ex_waddr,
    output io_ctrl_mem_rs1_ra,
    output[4:0] io_ctrl_mem_waddr,
    output[4:0] io_ctrl_wb_waddr,
    output[7:0] io_ctrl_status_ip,
    output[7:0] io_ctrl_status_im,
    output[6:0] io_ctrl_status_zero,
    output io_ctrl_status_er,
    output io_ctrl_status_vm,
    output io_ctrl_status_s64,
    output io_ctrl_status_u64,
    output io_ctrl_status_ef,
    output io_ctrl_status_pei,
    output io_ctrl_status_ei,
    output io_ctrl_status_ps,
    output io_ctrl_status_s,
    output io_ctrl_fp_sboard_clr,
    output[4:0] io_ctrl_fp_sboard_clra,
    output io_ctrl_csr_replay,
    input  io_dmem_req_ready,
    //output io_dmem_req_valid
    //output io_dmem_req_bits_kill
    //output[2:0] io_dmem_req_bits_typ
    //output io_dmem_req_bits_phys
    output[43:0] io_dmem_req_bits_addr,
    output[63:0] io_dmem_req_bits_data,
    output[7:0] io_dmem_req_bits_tag,
    //output[4:0] io_dmem_req_bits_cmd
    input  io_dmem_resp_valid,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [2:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [7:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_sret,
    output[7:0] io_ptw_status_ip,
    output[7:0] io_ptw_status_im,
    output[6:0] io_ptw_status_zero,
    output io_ptw_status_er,
    output io_ptw_status_vm,
    output io_ptw_status_s64,
    output io_ptw_status_u64,
    output io_ptw_status_ef,
    output io_ptw_status_pei,
    output io_ptw_status_ei,
    output io_ptw_status_ps,
    output io_ptw_status_s,
    //output io_imem_req_valid
    output[43:0] io_imem_req_bits_pc,
    //output io_imem_resp_ready
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input [42:0] io_imem_btb_resp_bits_target,
    input [2:0] io_imem_btb_resp_bits_entry,
    input [3:0] io_imem_btb_resp_bits_bht_index,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    //output io_imem_btb_update_valid
    //output io_imem_btb_update_bits_prediction_valid
    //output io_imem_btb_update_bits_prediction_bits_taken
    //output[42:0] io_imem_btb_update_bits_prediction_bits_target
    //output[2:0] io_imem_btb_update_bits_prediction_bits_entry
    //output[3:0] io_imem_btb_update_bits_prediction_bits_bht_index
    //output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value
    output[42:0] io_imem_btb_update_bits_pc,
    output[42:0] io_imem_btb_update_bits_target,
    output[42:0] io_imem_btb_update_bits_returnAddr,
    //output io_imem_btb_update_bits_taken
    //output io_imem_btb_update_bits_isJump
    //output io_imem_btb_update_bits_isCall
    //output io_imem_btb_update_bits_isReturn
    //output io_imem_btb_update_bits_incorrectTarget
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    //output io_imem_invalidate
    output[31:0] io_fpu_inst,
    output[63:0] io_fpu_fromint_data,
    output[2:0] io_fpu_fcsr_rm,
    input  io_fpu_fcsr_flags_valid,
    input [4:0] io_fpu_fcsr_flags_bits,
    input [63:0] io_fpu_store_data,
    input [63:0] io_fpu_toint_data,
    output io_fpu_dmem_resp_val,
    output[2:0] io_fpu_dmem_resp_type,
    output[4:0] io_fpu_dmem_resp_tag,
    output[63:0] io_fpu_dmem_resp_data,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[3:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [3:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    //output io_rocc_exception
);

  wire T0;
  wire[31:0] T1;
  reg [31:0] wb_reg_inst;
  wire[31:0] T2;
  reg [31:0] mem_reg_inst;
  wire[31:0] T3;
  reg [31:0] ex_reg_inst;
  wire[31:0] T4;
  wire T5;
  wire T6;
  reg  ex_reg_kill;
  wire T7;
  reg  mem_reg_kill;
  wire[31:0] T8;
  wire[63:0] T9;
  reg [63:0] R10;
  reg [63:0] R11;
  wire[63:0] ex_rs_1;
  wire[63:0] T12;
  reg [1:0] ex_reg_rs_lsb_1;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire[63:0] id_rs_1;
  wire[63:0] T16;
  wire[63:0] T17;
  reg [63:0] T18 [30:0];
  wire[63:0] T19;
  wire[63:0] wb_wdata;
  wire[63:0] T20;
  wire[63:0] T21;
  wire[63:0] T22;
  reg [63:0] wb_reg_wdata;
  wire[63:0] T23;
  wire[63:0] T24;
  wire[63:0] mem_int_wdata;
  reg [63:0] mem_reg_wdata;
  wire[63:0] T25;
  wire[63:0] alu_io_out;
  wire[63:0] T26;
  wire[44:0] mem_br_target;
  wire[44:0] T27;
  wire[44:0] T28;
  reg [43:0] mem_reg_pc;
  wire[43:0] T29;
  reg [43:0] ex_reg_pc;
  wire[43:0] T30;
  wire[44:0] T31;
  wire[21:0] T32;
  wire[21:0] T33;
  wire[21:0] T34;
  wire[21:0] T35;
  wire[11:0] T36;
  wire[4:0] T37;
  wire[3:0] T38;
  wire[6:0] T39;
  wire[5:0] T40;
  wire T41;
  wire T42;
  wire[9:0] T43;
  wire[8:0] T44;
  wire[7:0] T45;
  wire[7:0] T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire[21:0] T52;
  wire[14:0] T53;
  wire[14:0] T54;
  wire[11:0] T55;
  wire[4:0] T56;
  wire[3:0] T57;
  wire[6:0] T58;
  wire[5:0] T59;
  wire T60;
  wire T61;
  wire[2:0] T62;
  wire[1:0] T63;
  wire T64;
  wire T65;
  wire[6:0] T66;
  wire T67;
  wire T68;
  wire[22:0] T69;
  wire T70;
  wire[18:0] T71;
  wire T72;
  wire T73;
  wire[63:0] pcr_io_rw_rdata;
  wire T74;
  wire[63:0] ll_wdata;
  wire[63:0] div_io_resp_bits_data;
  wire T75;
  wire dmem_resp_xpu;
  wire T76;
  wire T77;
  wire dmem_resp_valid;
  wire T78;
  wire T79;
  wire[4:0] T80;
  wire[4:0] T81;
  wire[4:0] wb_waddr;
  wire T82;
  wire T83;
  wire wb_wen;
  wire[4:0] T84;
  wire[4:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg [61:0] ex_reg_rs_msb_1;
  wire[61:0] T90;
  wire[61:0] T91;
  wire T92;
  wire T93;
  wire[63:0] T94;
  wire[63:0] T95;
  wire[63:0] T96;
  wire bypass_0;
  wire[63:0] bypass_1;
  wire T97;
  wire[1:0] T98;
  wire[63:0] T99;
  wire[63:0] bypass_2;
  wire[63:0] bypass_3;
  wire T100;
  wire T101;
  reg  ex_reg_rs_bypass_1;
  wire T102;
  wire[4:0] T103;
  wire[4:0] T104;
  wire[63:0] T105;
  reg [63:0] R106;
  reg [63:0] R107;
  wire[63:0] ex_rs_0;
  wire[63:0] T108;
  reg [1:0] ex_reg_rs_lsb_0;
  wire[1:0] T109;
  wire[1:0] T110;
  wire[1:0] T111;
  wire[63:0] id_rs_0;
  wire[63:0] T112;
  wire[63:0] T113;
  wire[4:0] T114;
  wire[4:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  reg [61:0] ex_reg_rs_msb_0;
  wire[61:0] T120;
  wire[61:0] T121;
  wire T122;
  wire T123;
  wire[63:0] T124;
  wire[63:0] T125;
  wire[63:0] T126;
  wire T127;
  wire[1:0] T128;
  wire[63:0] T129;
  wire T130;
  wire T131;
  reg  ex_reg_rs_bypass_0;
  wire T132;
  wire[4:0] T133;
  wire[4:0] T134;
  wire T135;
  wire[63:0] T136;
  wire[4:0] T137;
  wire[4:0] T138;
  wire[43:0] T139;
  reg [43:0] wb_reg_pc;
  wire[43:0] T140;
  wire T141;
  wire[32:0] T142;
  wire[32:0] T143;
  wire[63:0] pcr_io_time;
  wire T144;
  wire[1135:0] T145;
  wire[63:0] T146;
  wire[63:0] T147;
  wire[63:0] T148;
  wire[63:0] T149;
  wire T150;
  wire[63:0] T151;
  wire T152;
  wire[1:0] T153;
  wire[11:0] T154;
  wire T155;
  wire T156;
  wire dmem_resp_replay;
  reg  ex_reg_ctrl_fn_dw;
  wire T157;
  wire T158;
  reg [3:0] ex_reg_ctrl_fn_alu;
  wire[3:0] T159;
  wire[63:0] ex_op1;
  wire[63:0] T160;
  wire[43:0] T161;
  wire[43:0] T162;
  wire T163;
  reg [1:0] ex_reg_sel_alu1;
  wire[1:0] T164;
  wire[19:0] T165;
  wire T166;
  wire[63:0] T167;
  wire T168;
  wire[63:0] T169;
  wire[63:0] ex_op2;
  wire[63:0] T170;
  wire[31:0] T171;
  wire[31:0] T172;
  wire[3:0] T173;
  wire T174;
  reg [2:0] ex_reg_sel_alu2;
  wire[2:0] T175;
  wire[27:0] T176;
  wire T177;
  wire[31:0] ex_imm;
  wire[31:0] T178;
  wire[11:0] T179;
  wire[4:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  reg [2:0] ex_reg_sel_imm;
  wire[2:0] T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire[3:0] T191;
  wire[3:0] T192;
  wire[3:0] T193;
  wire[3:0] T194;
  wire[3:0] T195;
  wire T196;
  wire[3:0] T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire[6:0] T202;
  wire[5:0] T203;
  wire[5:0] T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire[19:0] T222;
  wire[18:0] T223;
  wire[7:0] T224;
  wire[7:0] T225;
  wire[7:0] T226;
  wire[7:0] T227;
  wire T228;
  wire T229;
  wire T230;
  wire[10:0] T231;
  wire[10:0] T232;
  wire[10:0] T233;
  wire[10:0] T234;
  wire T235;
  wire T236;
  wire[31:0] T237;
  wire T238;
  wire[63:0] T239;
  wire T240;
  reg [63:0] wb_reg_rs2;
  wire[63:0] T241;
  reg [63:0] mem_reg_rs2;
  wire[63:0] T242;
  wire[6:0] T243;
  wire[4:0] T244;
  wire T245;
  wire T246;
  wire T247;
  wire[4:0] T248;
  wire[4:0] T249;
  wire[6:0] T250;
  wire[4:0] T251;
  wire[6:0] dmem_resp_waddr;
  wire[7:0] T252;
  wire T253;
  wire dmem_resp_fpu;
  wire T254;
  wire[2:0] pcr_io_fcsr_rm;
  wire[42:0] T255;
  wire[42:0] T256;
  wire[42:0] T257;
  wire[43:0] T258;
  wire[44:0] T259;
  wire[44:0] T260;
  wire[44:0] T261;
  wire[43:0] T262;
  wire[43:0] pcr_io_evec;
  wire T263;
  wire[44:0] mem_npc;
  wire[44:0] T264;
  wire[43:0] T265;
  wire[42:0] T266;
  wire T267;
  wire T268;
  wire T269;
  wire[1:0] T270;
  wire T271;
  wire T272;
  wire T273;
  wire[21:0] T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire pcr_io_status_s;
  wire pcr_io_status_ps;
  wire pcr_io_status_ei;
  wire pcr_io_status_pei;
  wire pcr_io_status_ef;
  wire pcr_io_status_u64;
  wire pcr_io_status_s64;
  wire pcr_io_status_vm;
  wire pcr_io_status_er;
  wire[6:0] pcr_io_status_zero;
  wire[7:0] pcr_io_status_im;
  wire[7:0] pcr_io_status_ip;
  wire pcr_io_fatc;
  wire[31:0] pcr_io_ptbr;
  wire[7:0] T281;
  wire[5:0] T282;
  wire[63:0] T283;
  wire[43:0] T284;
  wire[43:0] T285;
  wire[42:0] T286;
  wire[63:0] alu_io_adder_out;
  wire T287;
  wire T288;
  wire T289;
  wire[1:0] T290;
  wire T291;
  wire T292;
  wire T293;
  wire[21:0] T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire pcr_io_replay;
  wire[4:0] T300;
  wire T301;
  wire[4:0] T302;
  wire[4:0] T303;
  wire T304;
  wire[4:0] T305;
  wire[4:0] T306;
  wire[4:0] T307;
  wire[6:0] T308;
  wire[6:0] T309;
  wire[4:0] div_io_resp_bits_tag;
  wire T310;
  wire T311;
  wire div_io_resp_valid;
  wire div_io_req_ready;
  wire T312;
  wire[44:0] T313;
  wire[43:0] T314;
  wire T315;
  wire pcr_io_host_debug_stats_pcr;
  wire pcr_io_host_ipi_rep_ready;
  wire pcr_io_host_ipi_req_bits;
  wire pcr_io_host_ipi_req_valid;
  wire[63:0] pcr_io_host_pcr_rep_bits;
  wire pcr_io_host_pcr_rep_valid;
  wire pcr_io_host_pcr_req_ready;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    wb_reg_inst = {1{$random}};
    mem_reg_inst = {1{$random}};
    ex_reg_inst = {1{$random}};
    ex_reg_kill = {1{$random}};
    mem_reg_kill = {1{$random}};
    R10 = {2{$random}};
    R11 = {2{$random}};
    ex_reg_rs_lsb_1 = {1{$random}};
    for (initvar = 0; initvar < 31; initvar = initvar+1)
      T18[initvar] = {2{$random}};
    wb_reg_wdata = {2{$random}};
    mem_reg_wdata = {2{$random}};
    mem_reg_pc = {2{$random}};
    ex_reg_pc = {2{$random}};
    ex_reg_rs_msb_1 = {2{$random}};
    ex_reg_rs_bypass_1 = {1{$random}};
    R106 = {2{$random}};
    R107 = {2{$random}};
    ex_reg_rs_lsb_0 = {1{$random}};
    ex_reg_rs_msb_0 = {2{$random}};
    ex_reg_rs_bypass_0 = {1{$random}};
    wb_reg_pc = {2{$random}};
    ex_reg_ctrl_fn_dw = {1{$random}};
    ex_reg_ctrl_fn_alu = {1{$random}};
    ex_reg_sel_alu1 = {1{$random}};
    ex_reg_sel_alu2 = {1{$random}};
    ex_reg_sel_imm = {1{$random}};
    wb_reg_rs2 = {2{$random}};
    mem_reg_rs2 = {2{$random}};
  end
`endif

  assign T0 = reset ^ 1'h1;
  assign T1 = wb_reg_inst;
  assign T2 = T7 ? mem_reg_inst : wb_reg_inst;
  assign T3 = T6 ? ex_reg_inst : mem_reg_inst;
  assign T4 = T5 ? io_imem_resp_bits_data : ex_reg_inst;
  assign T5 = io_ctrl_killd ^ 1'h1;
  assign T6 = ex_reg_kill ^ 1'h1;
  assign T7 = mem_reg_kill ^ 1'h1;
  assign T8 = wb_reg_inst;
  assign T9 = R10;
  assign ex_rs_1 = ex_reg_rs_bypass_1 ? T94 : T12;
  assign T12 = {ex_reg_rs_msb_1, ex_reg_rs_lsb_1};
  assign T13 = T89 ? io_ctrl_bypass_src_1 : T14;
  assign T14 = T88 ? T15 : ex_reg_rs_lsb_1;
  assign T15 = id_rs_1[1'h1:1'h0];
  assign id_rs_1 = T16;
  assign T16 = T86 ? wb_wdata : T17;
  assign T17 = T18[T84];
  always @(posedge clk)
    if (T78)
      T18[T81] <= wb_wdata;
  assign wb_wdata = T20;
  assign T20 = T75 ? io_dmem_resp_bits_data_subword : T21;
  assign T21 = io_ctrl_ll_wen ? ll_wdata : T22;
  assign T22 = T74 ? pcr_io_rw_rdata : wb_reg_wdata;
  assign T23 = T7 ? T24 : wb_reg_wdata;
  assign T24 = T73 ? io_fpu_toint_data : mem_int_wdata;
  assign mem_int_wdata = io_ctrl_mem_jalr ? T26 : mem_reg_wdata;
  assign T25 = T6 ? alu_io_out : mem_reg_wdata;
  assign T26 = {T71, mem_br_target};
  assign mem_br_target = T31 + T27;
  assign T27 = T28;
  assign T28 = {1'h0, mem_reg_pc};
  assign T29 = T6 ? ex_reg_pc : mem_reg_pc;
  assign T30 = T5 ? io_imem_resp_bits_pc : ex_reg_pc;
  assign T31 = {T69, T32};
  assign T32 = T68 ? T52 : T33;
  assign T33 = T49 ? T34 : 22'h4;
  assign T34 = T35;
  assign T35 = {T43, T36};
  assign T36 = {T39, T37};
  assign T37 = {T38, 1'h0};
  assign T38 = mem_reg_inst[5'h18:5'h15];
  assign T39 = {T41, T40};
  assign T40 = mem_reg_inst[5'h1e:5'h19];
  assign T41 = T42;
  assign T42 = mem_reg_inst[5'h14:5'h14];
  assign T43 = {T47, T44};
  assign T44 = {T47, T45};
  assign T45 = T46;
  assign T46 = mem_reg_inst[5'h13:4'hc];
  assign T47 = T48;
  assign T48 = mem_reg_inst[5'h1f:5'h1f];
  assign T49 = T51 & T50;
  assign T50 = io_ctrl_mem_branch ^ 1'h1;
  assign T51 = io_ctrl_mem_jalr ^ 1'h1;
  assign T52 = {T66, T53};
  assign T53 = T54;
  assign T54 = {T62, T55};
  assign T55 = {T58, T56};
  assign T56 = {T57, 1'h0};
  assign T57 = mem_reg_inst[4'hb:4'h8];
  assign T58 = {T60, T59};
  assign T59 = mem_reg_inst[5'h1e:5'h19];
  assign T60 = T61;
  assign T61 = mem_reg_inst[3'h7:3'h7];
  assign T62 = {T64, T63};
  assign T63 = {T64, T64};
  assign T64 = T65;
  assign T65 = mem_reg_inst[5'h1f:5'h1f];
  assign T66 = T67 ? 7'h7f : 7'h0;
  assign T67 = T53[4'he:4'he];
  assign T68 = io_ctrl_mem_branch & io_ctrl_mem_br_taken;
  assign T69 = T70 ? 23'h7fffff : 23'h0;
  assign T70 = T32[5'h15:5'h15];
  assign T71 = T72 ? 19'h7ffff : 19'h0;
  assign T72 = mem_br_target[6'h2c:6'h2c];
  assign T73 = io_ctrl_mem_fp_val & io_ctrl_mem_wen;
  assign T74 = io_ctrl_csr != 3'h0;
  assign ll_wdata = div_io_resp_bits_data;
  assign T75 = dmem_resp_valid & dmem_resp_xpu;
  assign dmem_resp_xpu = T76 ^ 1'h1;
  assign T76 = T77;
  assign T77 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign T78 = T82 & T79;
  assign T79 = T80 < 5'h1f;
  assign T80 = T81[3'h4:1'h0];
  assign T81 = ~ wb_waddr;
  assign wb_waddr = io_ctrl_ll_wen ? io_ctrl_ll_waddr : io_ctrl_wb_waddr;
  assign T82 = wb_wen & T83;
  assign T83 = wb_waddr != 5'h0;
  assign wb_wen = io_ctrl_ll_wen | io_ctrl_wb_wen;
  assign T84 = ~ T85;
  assign T85 = io_imem_resp_bits_data[5'h18:5'h14];
  assign T86 = T82 & T87;
  assign T87 = wb_waddr == T85;
  assign T88 = T5 & io_ctrl_ren_1;
  assign T89 = T5 & io_ctrl_bypass_1;
  assign T90 = T92 ? T91 : ex_reg_rs_msb_1;
  assign T91 = id_rs_1 >> 2'h2;
  assign T92 = T88 & T93;
  assign T93 = io_ctrl_bypass_1 ^ 1'h1;
  assign T94 = T101 ? T99 : T95;
  assign T95 = T97 ? bypass_1 : T96;
  assign T96 = {63'h0, bypass_0};
  assign bypass_0 = 1'h0;
  assign bypass_1 = mem_reg_wdata;
  assign T97 = T98[1'h0:1'h0];
  assign T98 = ex_reg_rs_lsb_1;
  assign T99 = T100 ? bypass_3 : bypass_2;
  assign bypass_2 = wb_reg_wdata;
  assign bypass_3 = io_dmem_resp_bits_data;
  assign T100 = T98[1'h0:1'h0];
  assign T101 = T98[1'h1:1'h1];
  assign T102 = T5 ? io_ctrl_bypass_1 : ex_reg_rs_bypass_1;
  assign T103 = T104;
  assign T104 = wb_reg_inst[5'h18:5'h14];
  assign T105 = R106;
  assign ex_rs_0 = ex_reg_rs_bypass_0 ? T124 : T108;
  assign T108 = {ex_reg_rs_msb_0, ex_reg_rs_lsb_0};
  assign T109 = T119 ? io_ctrl_bypass_src_0 : T110;
  assign T110 = T118 ? T111 : ex_reg_rs_lsb_0;
  assign T111 = id_rs_0[1'h1:1'h0];
  assign id_rs_0 = T112;
  assign T112 = T116 ? wb_wdata : T113;
  assign T113 = T18[T114];
  assign T114 = ~ T115;
  assign T115 = io_imem_resp_bits_data[5'h13:4'hf];
  assign T116 = T82 & T117;
  assign T117 = wb_waddr == T115;
  assign T118 = T5 & io_ctrl_ren_0;
  assign T119 = T5 & io_ctrl_bypass_0;
  assign T120 = T122 ? T121 : ex_reg_rs_msb_0;
  assign T121 = id_rs_0 >> 2'h2;
  assign T122 = T118 & T123;
  assign T123 = io_ctrl_bypass_0 ^ 1'h1;
  assign T124 = T131 ? T129 : T125;
  assign T125 = T127 ? bypass_1 : T126;
  assign T126 = {63'h0, bypass_0};
  assign T127 = T128[1'h0:1'h0];
  assign T128 = ex_reg_rs_lsb_0;
  assign T129 = T130 ? bypass_3 : bypass_2;
  assign T130 = T128[1'h0:1'h0];
  assign T131 = T128[1'h1:1'h1];
  assign T132 = T5 ? io_ctrl_bypass_0 : ex_reg_rs_bypass_0;
  assign T133 = T134;
  assign T134 = wb_reg_inst[5'h13:4'hf];
  assign T135 = wb_wen;
  assign T136 = wb_wdata;
  assign T137 = T138;
  assign T138 = wb_wen ? wb_waddr : 5'h0;
  assign T139 = wb_reg_pc;
  assign T140 = T7 ? mem_reg_pc : wb_reg_pc;
  assign T141 = io_ctrl_retire;
  assign T142 = T143;
  assign T143 = pcr_io_time[6'h20:1'h0];
  assign T144 = io_host_id;
  assign T146 = T152 ? T151 : T147;
  assign T147 = T150 ? T148 : wb_reg_wdata;
  assign T148 = pcr_io_rw_rdata & T149;
  assign T149 = ~ wb_reg_wdata;
  assign T150 = io_ctrl_csr == 3'h3;
  assign T151 = pcr_io_rw_rdata | wb_reg_wdata;
  assign T152 = io_ctrl_csr == 3'h2;
  assign T153 = io_ctrl_csr[1'h1:1'h0];
  assign T154 = wb_reg_inst[5'h1f:5'h14];
  assign T155 = T156 ? 1'h0 : io_ctrl_ll_ready;
  assign T156 = dmem_resp_replay & dmem_resp_xpu;
  assign dmem_resp_replay = io_dmem_resp_bits_replay & io_dmem_resp_bits_has_data;
  assign T157 = T5 ? T158 : ex_reg_ctrl_fn_dw;
  assign T158 = io_ctrl_fn_dw;
  assign T159 = T5 ? io_ctrl_fn_alu : ex_reg_ctrl_fn_alu;
  assign ex_op1 = T168 ? T167 : T160;
  assign T160 = {T165, T161};
  assign T161 = T163 ? T162 : 44'h0;
  assign T162 = ex_reg_pc;
  assign T163 = ex_reg_sel_alu1 == 2'h2;
  assign T164 = T5 ? io_ctrl_sel_alu1 : ex_reg_sel_alu1;
  assign T165 = T166 ? 20'hfffff : 20'h0;
  assign T166 = T161[6'h2b:6'h2b];
  assign T167 = ex_rs_0;
  assign T168 = ex_reg_sel_alu1 == 2'h1;
  assign T169 = ex_op2;
  assign ex_op2 = T240 ? T239 : T170;
  assign T170 = {T237, T171};
  assign T171 = T236 ? ex_imm : T172;
  assign T172 = {T176, T173};
  assign T173 = T174 ? 4'h4 : 4'h0;
  assign T174 = ex_reg_sel_alu2 == 3'h1;
  assign T175 = T5 ? io_ctrl_sel_alu2 : ex_reg_sel_alu2;
  assign T176 = T177 ? 28'hfffffff : 28'h0;
  assign T177 = T173[2'h3:2'h3];
  assign ex_imm = T178;
  assign T178 = {T222, T179};
  assign T179 = {T202, T180};
  assign T180 = {T191, T181};
  assign T181 = T190 ? T189 : T182;
  assign T182 = T188 ? T187 : T183;
  assign T183 = T185 ? T184 : 1'h0;
  assign T184 = ex_reg_inst[4'hf:4'hf];
  assign T185 = ex_reg_sel_imm == 3'h5;
  assign T186 = T5 ? io_ctrl_sel_imm : ex_reg_sel_imm;
  assign T187 = ex_reg_inst[5'h14:5'h14];
  assign T188 = ex_reg_sel_imm == 3'h4;
  assign T189 = ex_reg_inst[3'h7:3'h7];
  assign T190 = ex_reg_sel_imm == 3'h0;
  assign T191 = T201 ? 4'h0 : T192;
  assign T192 = T198 ? T197 : T193;
  assign T193 = T196 ? T195 : T194;
  assign T194 = ex_reg_inst[5'h18:5'h15];
  assign T195 = ex_reg_inst[5'h13:5'h10];
  assign T196 = ex_reg_sel_imm == 3'h5;
  assign T197 = ex_reg_inst[4'hb:4'h8];
  assign T198 = T200 | T199;
  assign T199 = ex_reg_sel_imm == 3'h1;
  assign T200 = ex_reg_sel_imm == 3'h0;
  assign T201 = ex_reg_sel_imm == 3'h2;
  assign T202 = {T208, T203};
  assign T203 = T205 ? 6'h0 : T204;
  assign T204 = ex_reg_inst[5'h1e:5'h19];
  assign T205 = T207 | T206;
  assign T206 = ex_reg_sel_imm == 3'h5;
  assign T207 = ex_reg_sel_imm == 3'h2;
  assign T208 = T219 ? 1'h0 : T209;
  assign T209 = T218 ? T216 : T210;
  assign T210 = T215 ? T213 : T211;
  assign T211 = T212;
  assign T212 = ex_reg_inst[5'h1f:5'h1f];
  assign T213 = T214;
  assign T214 = ex_reg_inst[3'h7:3'h7];
  assign T215 = ex_reg_sel_imm == 3'h1;
  assign T216 = T217;
  assign T217 = ex_reg_inst[5'h14:5'h14];
  assign T218 = ex_reg_sel_imm == 3'h3;
  assign T219 = T221 | T220;
  assign T220 = ex_reg_sel_imm == 3'h5;
  assign T221 = ex_reg_sel_imm == 3'h2;
  assign T222 = {T211, T223};
  assign T223 = {T231, T224};
  assign T224 = T228 ? T227 : T225;
  assign T225 = T226;
  assign T226 = ex_reg_inst[5'h13:4'hc];
  assign T227 = T211 ? 8'hff : 8'h0;
  assign T228 = T230 & T229;
  assign T229 = ex_reg_sel_imm != 3'h3;
  assign T230 = ex_reg_sel_imm != 3'h2;
  assign T231 = T235 ? T233 : T232;
  assign T232 = T211 ? 11'h7ff : 11'h0;
  assign T233 = T234;
  assign T234 = ex_reg_inst[5'h1e:5'h14];
  assign T235 = ex_reg_sel_imm == 3'h2;
  assign T236 = ex_reg_sel_alu2 == 3'h3;
  assign T237 = T238 ? 32'hffffffff : 32'h0;
  assign T238 = T171[5'h1f:5'h1f];
  assign T239 = ex_rs_1;
  assign T240 = ex_reg_sel_alu2 == 3'h2;
  assign io_rocc_cmd_bits_rs2 = wb_reg_rs2;
  assign T241 = io_ctrl_mem_rocc_val ? mem_reg_rs2 : wb_reg_rs2;
  assign T242 = io_ctrl_ex_rs2_val ? ex_rs_1 : mem_reg_rs2;
  assign io_rocc_cmd_bits_rs1 = wb_reg_wdata;
  assign io_rocc_cmd_bits_inst_opcode = T243;
  assign T243 = wb_reg_inst[3'h6:1'h0];
  assign io_rocc_cmd_bits_inst_rd = T244;
  assign T244 = wb_reg_inst[4'hb:3'h7];
  assign io_rocc_cmd_bits_inst_xs2 = T245;
  assign T245 = wb_reg_inst[4'hc:4'hc];
  assign io_rocc_cmd_bits_inst_xs1 = T246;
  assign T246 = wb_reg_inst[4'hd:4'hd];
  assign io_rocc_cmd_bits_inst_xd = T247;
  assign T247 = wb_reg_inst[4'he:4'he];
  assign io_rocc_cmd_bits_inst_rs1 = T248;
  assign T248 = wb_reg_inst[5'h13:4'hf];
  assign io_rocc_cmd_bits_inst_rs2 = T249;
  assign T249 = wb_reg_inst[5'h18:5'h14];
  assign io_rocc_cmd_bits_inst_funct = T250;
  assign T250 = wb_reg_inst[5'h1f:5'h19];
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data;
  assign io_fpu_dmem_resp_tag = T251;
  assign T251 = dmem_resp_waddr[3'h4:1'h0];
  assign dmem_resp_waddr = T252 >> 1'h1;
  assign T252 = io_dmem_resp_bits_tag;
  assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ;
  assign io_fpu_dmem_resp_val = T253;
  assign T253 = dmem_resp_valid & dmem_resp_fpu;
  assign dmem_resp_fpu = T254;
  assign T254 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign io_fpu_fcsr_rm = pcr_io_fcsr_rm;
  assign io_fpu_fromint_data = ex_rs_0;
  assign io_fpu_inst = io_imem_resp_bits_data;
  assign io_imem_btb_update_bits_returnAddr = T255;
  assign T255 = mem_int_wdata[6'h2a:1'h0];
  assign io_imem_btb_update_bits_target = T256;
  assign T256 = io_imem_req_bits_pc[6'h2a:1'h0];
  assign io_imem_btb_update_bits_pc = T257;
  assign T257 = mem_reg_pc[6'h2a:1'h0];
  assign io_imem_req_bits_pc = T258;
  assign T258 = T259[6'h2b:1'h0];
  assign T259 = T260;
  assign T260 = T280 ? mem_npc : T261;
  assign T261 = {1'h0, T262};
  assign T262 = T263 ? pcr_io_evec : wb_reg_pc;
  assign T263 = io_ctrl_sel_pc == 3'h3;
  assign mem_npc = io_ctrl_mem_jalr ? T264 : mem_br_target;
  assign T264 = {1'h0, T265};
  assign T265 = {T267, T266};
  assign T266 = mem_reg_wdata[6'h2a:1'h0];
  assign T267 = T277 ? T276 : T268;
  assign T268 = T272 ? T271 : T269;
  assign T269 = T270[1'h0:1'h0];
  assign T270 = mem_reg_wdata[6'h2b:6'h2a];
  assign T271 = T270 == 2'h3;
  assign T272 = T275 | T273;
  assign T273 = T274 == 22'h3ffffe;
  assign T274 = mem_reg_wdata >> 6'h2a;
  assign T275 = T274 == 22'h3fffff;
  assign T276 = T270 != 2'h0;
  assign T277 = T279 | T278;
  assign T278 = T274 == 22'h1;
  assign T279 = T274 == 22'h0;
  assign T280 = io_ctrl_sel_pc == 3'h1;
  assign io_ptw_status_s = pcr_io_status_s;
  assign io_ptw_status_ps = pcr_io_status_ps;
  assign io_ptw_status_ei = pcr_io_status_ei;
  assign io_ptw_status_pei = pcr_io_status_pei;
  assign io_ptw_status_ef = pcr_io_status_ef;
  assign io_ptw_status_u64 = pcr_io_status_u64;
  assign io_ptw_status_s64 = pcr_io_status_s64;
  assign io_ptw_status_vm = pcr_io_status_vm;
  assign io_ptw_status_er = pcr_io_status_er;
  assign io_ptw_status_zero = pcr_io_status_zero;
  assign io_ptw_status_im = pcr_io_status_im;
  assign io_ptw_status_ip = pcr_io_status_ip;
  assign io_ptw_sret = io_ctrl_sret;
  assign io_ptw_invalidate = pcr_io_fatc;
  assign io_ptw_ptbr = pcr_io_ptbr;
  assign io_dmem_req_bits_tag = T281;
  assign T281 = {2'h0, T282};
  assign T282 = {io_ctrl_ex_waddr, io_ctrl_ex_fp_val};
  assign io_dmem_req_bits_data = T283;
  assign T283 = io_ctrl_mem_fp_val ? io_fpu_store_data : mem_reg_rs2;
  assign io_dmem_req_bits_addr = T284;
  assign T284 = T285;
  assign T285 = {T287, T286};
  assign T286 = alu_io_adder_out[6'h2a:1'h0];
  assign T287 = T297 ? T296 : T288;
  assign T288 = T292 ? T291 : T289;
  assign T289 = T290[1'h0:1'h0];
  assign T290 = alu_io_adder_out[6'h2b:6'h2a];
  assign T291 = T290 == 2'h3;
  assign T292 = T295 | T293;
  assign T293 = T294 == 22'h3ffffe;
  assign T294 = ex_rs_0 >> 6'h2a;
  assign T295 = T294 == 22'h3fffff;
  assign T296 = T290 != 2'h0;
  assign T297 = T299 | T298;
  assign T298 = T294 == 22'h1;
  assign T299 = T294 == 22'h0;
  assign io_ctrl_csr_replay = pcr_io_replay;
  assign io_ctrl_fp_sboard_clra = T300;
  assign T300 = dmem_resp_waddr[3'h4:1'h0];
  assign io_ctrl_fp_sboard_clr = T301;
  assign T301 = dmem_resp_replay & dmem_resp_fpu;
  assign io_ctrl_status_s = pcr_io_status_s;
  assign io_ctrl_status_ps = pcr_io_status_ps;
  assign io_ctrl_status_ei = pcr_io_status_ei;
  assign io_ctrl_status_pei = pcr_io_status_pei;
  assign io_ctrl_status_ef = pcr_io_status_ef;
  assign io_ctrl_status_u64 = pcr_io_status_u64;
  assign io_ctrl_status_s64 = pcr_io_status_s64;
  assign io_ctrl_status_vm = pcr_io_status_vm;
  assign io_ctrl_status_er = pcr_io_status_er;
  assign io_ctrl_status_zero = pcr_io_status_zero;
  assign io_ctrl_status_im = pcr_io_status_im;
  assign io_ctrl_status_ip = pcr_io_status_ip;
  assign io_ctrl_wb_waddr = T302;
  assign T302 = wb_reg_inst[4'hb:3'h7];
  assign io_ctrl_mem_waddr = T303;
  assign T303 = mem_reg_inst[4'hb:3'h7];
  assign io_ctrl_mem_rs1_ra = T304;
  assign T304 = T305 == 5'h1;
  assign T305 = mem_reg_inst[5'h13:4'hf];
  assign io_ctrl_ex_waddr = T306;
  assign T306 = ex_reg_inst[4'hb:3'h7];
  assign io_ctrl_ll_waddr = T307;
  assign T307 = T308[3'h4:1'h0];
  assign T308 = T156 ? dmem_resp_waddr : T309;
  assign T309 = {2'h0, div_io_resp_bits_tag};
  assign io_ctrl_ll_wen = T310;
  assign T310 = T156 ? 1'h1 : T311;
  assign T311 = T155 & div_io_resp_valid;
  assign io_ctrl_div_mul_rdy = div_io_req_ready;
  assign io_ctrl_mem_misprediction = T312;
  assign T312 = mem_npc != T313;
  assign T313 = {1'h0, T314};
  assign T314 = io_ctrl_ex_valid ? ex_reg_pc : io_imem_resp_bits_pc;
  assign io_ctrl_mem_br_taken = T315;
  assign T315 = mem_reg_wdata[1'h0:1'h0];
  assign io_ctrl_inst = io_imem_resp_bits_data;
  assign io_host_debug_stats_pcr = pcr_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = pcr_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = pcr_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = pcr_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = pcr_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = pcr_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = pcr_io_host_pcr_req_ready;
  ALU alu(
       .io_dw( ex_reg_ctrl_fn_dw ),
       .io_fn( ex_reg_ctrl_fn_alu ),
       .io_in2( T169 ),
       .io_in1( ex_op1 ),
       .io_out( alu_io_out ),
       .io_adder_out( alu_io_adder_out )
  );
  MulDiv div(.clk(clk), .reset(reset),
       .io_req_ready( div_io_req_ready ),
       .io_req_valid( io_ctrl_div_mul_val ),
       .io_req_bits_fn( ex_reg_ctrl_fn_alu ),
       .io_req_bits_dw( ex_reg_ctrl_fn_dw ),
       .io_req_bits_in1( ex_rs_0 ),
       .io_req_bits_in2( ex_rs_1 ),
       .io_req_bits_tag( io_ctrl_ex_waddr ),
       .io_kill( io_ctrl_div_mul_kill ),
       .io_resp_ready( T155 ),
       .io_resp_valid( div_io_resp_valid ),
       .io_resp_bits_data( div_io_resp_bits_data ),
       .io_resp_bits_tag( div_io_resp_bits_tag )
  );
  CSRFile pcr(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( pcr_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( pcr_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( pcr_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( pcr_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( pcr_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( pcr_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( pcr_io_host_debug_stats_pcr ),
       .io_rw_addr( T154 ),
       .io_rw_cmd( T153 ),
       .io_rw_rdata( pcr_io_rw_rdata ),
       .io_rw_wdata( T146 ),
       .io_status_ip( pcr_io_status_ip ),
       .io_status_im( pcr_io_status_im ),
       .io_status_zero( pcr_io_status_zero ),
       .io_status_er( pcr_io_status_er ),
       .io_status_vm( pcr_io_status_vm ),
       .io_status_s64( pcr_io_status_s64 ),
       .io_status_u64( pcr_io_status_u64 ),
       .io_status_ef( pcr_io_status_ef ),
       .io_status_pei( pcr_io_status_pei ),
       .io_status_ei( pcr_io_status_ei ),
       .io_status_ps( pcr_io_status_ps ),
       .io_status_s( pcr_io_status_s ),
       .io_ptbr( pcr_io_ptbr ),
       .io_evec( pcr_io_evec ),
       .io_exception( io_ctrl_exception ),
       .io_retire( io_ctrl_retire ),
       .io_cause( io_ctrl_cause ),
       .io_badvaddr_wen( io_ctrl_badvaddr_wen ),
       .io_pc( wb_reg_pc ),
       .io_sret( io_ctrl_sret ),
       .io_fatc( pcr_io_fatc ),
       .io_replay( pcr_io_replay ),
       .io_time( pcr_io_time ),
       .io_fcsr_rm( pcr_io_fcsr_rm ),
       .io_fcsr_flags_valid( io_fpu_fcsr_flags_valid ),
       .io_fcsr_flags_bits( io_fpu_fcsr_flags_bits ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_write_mask( io_rocc_imem_acquire_bits_payload_write_mask ),
       .io_rocc_imem_acquire_bits_payload_subword_addr( io_rocc_imem_acquire_bits_payload_subword_addr ),
       .io_rocc_imem_acquire_bits_payload_atomic_opcode( io_rocc_imem_acquire_bits_payload_atomic_opcode ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
  );

  always @(posedge clk) begin
    if(T7) begin
      wb_reg_inst <= mem_reg_inst;
    end
    if(T6) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if(T5) begin
      ex_reg_inst <= io_imem_resp_bits_data;
    end
    ex_reg_kill <= io_ctrl_killd;
    mem_reg_kill <= ex_reg_kill;
    R10 <= R11;
    if(ex_reg_rs_bypass_1) begin
      R11 <= T94;
    end else begin
      R11 <= T12;
    end
    if(T89) begin
      ex_reg_rs_lsb_1 <= io_ctrl_bypass_src_1;
    end else if(T88) begin
      ex_reg_rs_lsb_1 <= T15;
    end
    if(T7) begin
      wb_reg_wdata <= T24;
    end
    if(T6) begin
      mem_reg_wdata <= alu_io_out;
    end
    if(T6) begin
      mem_reg_pc <= ex_reg_pc;
    end
    if(T5) begin
      ex_reg_pc <= io_imem_resp_bits_pc;
    end
    if(T92) begin
      ex_reg_rs_msb_1 <= T91;
    end
    if(T5) begin
      ex_reg_rs_bypass_1 <= io_ctrl_bypass_1;
    end
    R106 <= R107;
    if(ex_reg_rs_bypass_0) begin
      R107 <= T124;
    end else begin
      R107 <= T108;
    end
    if(T119) begin
      ex_reg_rs_lsb_0 <= io_ctrl_bypass_src_0;
    end else if(T118) begin
      ex_reg_rs_lsb_0 <= T111;
    end
    if(T122) begin
      ex_reg_rs_msb_0 <= T121;
    end
    if(T5) begin
      ex_reg_rs_bypass_0 <= io_ctrl_bypass_0;
    end
    if(T7) begin
      wb_reg_pc <= mem_reg_pc;
    end
    if(T5) begin
      ex_reg_ctrl_fn_dw <= T158;
    end
    if(T5) begin
      ex_reg_ctrl_fn_alu <= io_ctrl_fn_alu;
    end
    if(T5) begin
      ex_reg_sel_alu1 <= io_ctrl_sel_alu1;
    end
    if(T5) begin
      ex_reg_sel_alu2 <= io_ctrl_sel_alu2;
    end
    if(T5) begin
      ex_reg_sel_imm <= io_ctrl_sel_imm;
    end
    if(io_ctrl_mem_rocc_val) begin
      wb_reg_rs2 <= mem_reg_rs2;
    end
    if(io_ctrl_ex_rs2_val) begin
      mem_reg_rs2 <= ex_rs_1;
    end
`ifndef SYNTHESIS
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T0)
        $fwrite(32'h80000002, "C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n", T144, T142, T141, T139, T137, T136, T135, T133, T105, T103, T9, T8, T1);
`endif
  end
endmodule

module Core(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    output io_imem_req_valid,
    output[43:0] io_imem_req_bits_pc,
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input [42:0] io_imem_btb_resp_bits_target,
    input [2:0] io_imem_btb_resp_bits_entry,
    input [3:0] io_imem_btb_resp_bits_bht_index,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output[42:0] io_imem_btb_update_bits_prediction_bits_target,
    output[2:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[3:0] io_imem_btb_update_bits_prediction_bits_bht_index,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    output[42:0] io_imem_btb_update_bits_pc,
    output[42:0] io_imem_btb_update_bits_target,
    output[42:0] io_imem_btb_update_bits_returnAddr,
    output io_imem_btb_update_bits_taken,
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isCall,
    output io_imem_btb_update_bits_isReturn,
    output io_imem_btb_update_bits_incorrectTarget,
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    output io_imem_invalidate,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output io_dmem_req_bits_kill,
    output[2:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_phys,
    output[43:0] io_dmem_req_bits_addr,
    output[63:0] io_dmem_req_bits_data,
    output[7:0] io_dmem_req_bits_tag,
    output[4:0] io_dmem_req_bits_cmd,
    input  io_dmem_resp_valid,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [2:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [7:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_sret,
    output[7:0] io_ptw_status_ip,
    output[7:0] io_ptw_status_im,
    output[6:0] io_ptw_status_zero,
    output io_ptw_status_er,
    output io_ptw_status_vm,
    output io_ptw_status_s64,
    output io_ptw_status_u64,
    output io_ptw_status_ef,
    output io_ptw_status_pei,
    output io_ptw_status_ei,
    output io_ptw_status_ps,
    output io_ptw_status_s,
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[3:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [3:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    output io_rocc_exception
);

  wire ctrl_io_dpath_badvaddr_wen;
  wire[63:0] ctrl_io_dpath_cause;
  wire ctrl_io_dpath_exception;
  wire ctrl_io_dpath_retire;
  wire ctrl_io_dpath_ll_ready;
  wire[1:0] ctrl_io_dpath_bypass_src_0;
  wire[1:0] ctrl_io_dpath_bypass_src_1;
  wire ctrl_io_dpath_bypass_0;
  wire ctrl_io_dpath_bypass_1;
  wire ctrl_io_dpath_mem_rocc_val;
  wire ctrl_io_dpath_ex_rocc_val;
  wire ctrl_io_dpath_ex_rs2_val;
  wire[2:0] ctrl_io_dpath_ex_mem_type;
  wire ctrl_io_dpath_wb_wen;
  wire ctrl_io_dpath_mem_wen;
  wire ctrl_io_dpath_mem_branch;
  wire ctrl_io_dpath_mem_jalr;
  wire ctrl_io_dpath_ex_valid;
  wire ctrl_io_dpath_ex_wen;
  wire ctrl_io_dpath_mem_fp_val;
  wire ctrl_io_dpath_ex_fp_val;
  wire ctrl_io_dpath_wb_load;
  wire ctrl_io_dpath_mem_load;
  wire ctrl_io_dpath_sret;
  wire[2:0] ctrl_io_dpath_csr;
  wire ctrl_io_dpath_div_mul_kill;
  wire ctrl_io_dpath_div_mul_val;
  wire[3:0] ctrl_io_dpath_fn_alu;
  wire ctrl_io_dpath_fn_dw;
  wire[2:0] ctrl_io_dpath_sel_imm;
  wire[1:0] ctrl_io_dpath_sel_alu1;
  wire[2:0] ctrl_io_dpath_sel_alu2;
  wire ctrl_io_dpath_ren_0;
  wire ctrl_io_dpath_ren_1;
  wire ctrl_io_dpath_killd;
  wire[2:0] ctrl_io_dpath_sel_pc;
  wire dpath_io_ctrl_csr_replay;
  wire[4:0] dpath_io_ctrl_fp_sboard_clra;
  wire dpath_io_ctrl_fp_sboard_clr;
  wire dpath_io_ctrl_status_s;
  wire dpath_io_ctrl_status_ps;
  wire dpath_io_ctrl_status_ei;
  wire dpath_io_ctrl_status_pei;
  wire dpath_io_ctrl_status_ef;
  wire dpath_io_ctrl_status_u64;
  wire dpath_io_ctrl_status_s64;
  wire dpath_io_ctrl_status_vm;
  wire dpath_io_ctrl_status_er;
  wire[6:0] dpath_io_ctrl_status_zero;
  wire[7:0] dpath_io_ctrl_status_im;
  wire[7:0] dpath_io_ctrl_status_ip;
  wire[4:0] dpath_io_ctrl_wb_waddr;
  wire[4:0] dpath_io_ctrl_mem_waddr;
  wire dpath_io_ctrl_mem_rs1_ra;
  wire[4:0] dpath_io_ctrl_ex_waddr;
  wire[4:0] dpath_io_ctrl_ll_waddr;
  wire dpath_io_ctrl_ll_wen;
  wire dpath_io_ctrl_div_mul_rdy;
  wire dpath_io_ctrl_mem_misprediction;
  wire dpath_io_ctrl_mem_br_taken;
  wire[31:0] dpath_io_ctrl_inst;
  wire ctrl_io_rocc_exception;
  wire ctrl_io_rocc_s;
  wire[63:0] dpath_io_rocc_cmd_bits_rs2;
  wire[63:0] dpath_io_rocc_cmd_bits_rs1;
  wire[6:0] dpath_io_rocc_cmd_bits_inst_opcode;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rd;
  wire dpath_io_rocc_cmd_bits_inst_xs2;
  wire dpath_io_rocc_cmd_bits_inst_xs1;
  wire dpath_io_rocc_cmd_bits_inst_xd;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rs1;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rs2;
  wire[6:0] dpath_io_rocc_cmd_bits_inst_funct;
  wire ctrl_io_rocc_cmd_valid;
  wire dpath_io_ptw_status_s;
  wire dpath_io_ptw_status_ps;
  wire dpath_io_ptw_status_ei;
  wire dpath_io_ptw_status_pei;
  wire dpath_io_ptw_status_ef;
  wire dpath_io_ptw_status_u64;
  wire dpath_io_ptw_status_s64;
  wire dpath_io_ptw_status_vm;
  wire dpath_io_ptw_status_er;
  wire[6:0] dpath_io_ptw_status_zero;
  wire[7:0] dpath_io_ptw_status_im;
  wire[7:0] dpath_io_ptw_status_ip;
  wire dpath_io_ptw_sret;
  wire dpath_io_ptw_invalidate;
  wire[31:0] dpath_io_ptw_ptbr;
  wire[4:0] ctrl_io_dmem_req_bits_cmd;
  wire[7:0] dpath_io_dmem_req_bits_tag;
  wire[63:0] dpath_io_dmem_req_bits_data;
  wire[43:0] dpath_io_dmem_req_bits_addr;
  wire ctrl_io_dmem_req_bits_phys;
  wire[2:0] ctrl_io_dmem_req_bits_typ;
  wire ctrl_io_dmem_req_bits_kill;
  wire ctrl_io_dmem_req_valid;
  wire ctrl_io_imem_invalidate;
  wire ctrl_io_imem_btb_update_bits_incorrectTarget;
  wire ctrl_io_imem_btb_update_bits_isReturn;
  wire ctrl_io_imem_btb_update_bits_isCall;
  wire ctrl_io_imem_btb_update_bits_isJump;
  wire ctrl_io_imem_btb_update_bits_taken;
  wire[42:0] dpath_io_imem_btb_update_bits_returnAddr;
  wire[42:0] dpath_io_imem_btb_update_bits_target;
  wire[42:0] dpath_io_imem_btb_update_bits_pc;
  wire[1:0] ctrl_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire[3:0] ctrl_io_imem_btb_update_bits_prediction_bits_bht_index;
  wire[2:0] ctrl_io_imem_btb_update_bits_prediction_bits_entry;
  wire[42:0] ctrl_io_imem_btb_update_bits_prediction_bits_target;
  wire ctrl_io_imem_btb_update_bits_prediction_bits_taken;
  wire ctrl_io_imem_btb_update_bits_prediction_valid;
  wire ctrl_io_imem_btb_update_valid;
  wire ctrl_io_imem_resp_ready;
  wire[43:0] dpath_io_imem_req_bits_pc;
  wire ctrl_io_imem_req_valid;
  wire dpath_io_host_debug_stats_pcr;
  wire dpath_io_host_ipi_rep_ready;
  wire dpath_io_host_ipi_req_bits;
  wire dpath_io_host_ipi_req_valid;
  wire[63:0] dpath_io_host_pcr_rep_bits;
  wire dpath_io_host_pcr_rep_valid;
  wire dpath_io_host_pcr_req_ready;


  assign io_rocc_exception = ctrl_io_rocc_exception;
  assign io_rocc_s = ctrl_io_rocc_s;
  assign io_rocc_cmd_bits_rs2 = dpath_io_rocc_cmd_bits_rs2;
  assign io_rocc_cmd_bits_rs1 = dpath_io_rocc_cmd_bits_rs1;
  assign io_rocc_cmd_bits_inst_opcode = dpath_io_rocc_cmd_bits_inst_opcode;
  assign io_rocc_cmd_bits_inst_rd = dpath_io_rocc_cmd_bits_inst_rd;
  assign io_rocc_cmd_bits_inst_xs2 = dpath_io_rocc_cmd_bits_inst_xs2;
  assign io_rocc_cmd_bits_inst_xs1 = dpath_io_rocc_cmd_bits_inst_xs1;
  assign io_rocc_cmd_bits_inst_xd = dpath_io_rocc_cmd_bits_inst_xd;
  assign io_rocc_cmd_bits_inst_rs1 = dpath_io_rocc_cmd_bits_inst_rs1;
  assign io_rocc_cmd_bits_inst_rs2 = dpath_io_rocc_cmd_bits_inst_rs2;
  assign io_rocc_cmd_bits_inst_funct = dpath_io_rocc_cmd_bits_inst_funct;
  assign io_rocc_cmd_valid = ctrl_io_rocc_cmd_valid;
  assign io_ptw_status_s = dpath_io_ptw_status_s;
  assign io_ptw_status_ps = dpath_io_ptw_status_ps;
  assign io_ptw_status_ei = dpath_io_ptw_status_ei;
  assign io_ptw_status_pei = dpath_io_ptw_status_pei;
  assign io_ptw_status_ef = dpath_io_ptw_status_ef;
  assign io_ptw_status_u64 = dpath_io_ptw_status_u64;
  assign io_ptw_status_s64 = dpath_io_ptw_status_s64;
  assign io_ptw_status_vm = dpath_io_ptw_status_vm;
  assign io_ptw_status_er = dpath_io_ptw_status_er;
  assign io_ptw_status_zero = dpath_io_ptw_status_zero;
  assign io_ptw_status_im = dpath_io_ptw_status_im;
  assign io_ptw_status_ip = dpath_io_ptw_status_ip;
  assign io_ptw_sret = dpath_io_ptw_sret;
  assign io_ptw_invalidate = dpath_io_ptw_invalidate;
  assign io_ptw_ptbr = dpath_io_ptw_ptbr;
  assign io_dmem_req_bits_cmd = ctrl_io_dmem_req_bits_cmd;
  assign io_dmem_req_bits_tag = dpath_io_dmem_req_bits_tag;
  assign io_dmem_req_bits_data = dpath_io_dmem_req_bits_data;
  assign io_dmem_req_bits_addr = dpath_io_dmem_req_bits_addr;
  assign io_dmem_req_bits_phys = ctrl_io_dmem_req_bits_phys;
  assign io_dmem_req_bits_typ = ctrl_io_dmem_req_bits_typ;
  assign io_dmem_req_bits_kill = ctrl_io_dmem_req_bits_kill;
  assign io_dmem_req_valid = ctrl_io_dmem_req_valid;
  assign io_imem_invalidate = ctrl_io_imem_invalidate;
  assign io_imem_btb_update_bits_incorrectTarget = ctrl_io_imem_btb_update_bits_incorrectTarget;
  assign io_imem_btb_update_bits_isReturn = ctrl_io_imem_btb_update_bits_isReturn;
  assign io_imem_btb_update_bits_isCall = ctrl_io_imem_btb_update_bits_isCall;
  assign io_imem_btb_update_bits_isJump = ctrl_io_imem_btb_update_bits_isJump;
  assign io_imem_btb_update_bits_taken = ctrl_io_imem_btb_update_bits_taken;
  assign io_imem_btb_update_bits_returnAddr = dpath_io_imem_btb_update_bits_returnAddr;
  assign io_imem_btb_update_bits_target = dpath_io_imem_btb_update_bits_target;
  assign io_imem_btb_update_bits_pc = dpath_io_imem_btb_update_bits_pc;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = ctrl_io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_btb_update_bits_prediction_bits_bht_index = ctrl_io_imem_btb_update_bits_prediction_bits_bht_index;
  assign io_imem_btb_update_bits_prediction_bits_entry = ctrl_io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = ctrl_io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_btb_update_bits_prediction_bits_taken = ctrl_io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_btb_update_bits_prediction_valid = ctrl_io_imem_btb_update_bits_prediction_valid;
  assign io_imem_btb_update_valid = ctrl_io_imem_btb_update_valid;
  assign io_imem_resp_ready = ctrl_io_imem_resp_ready;
  assign io_imem_req_bits_pc = dpath_io_imem_req_bits_pc;
  assign io_imem_req_valid = ctrl_io_imem_req_valid;
  assign io_host_debug_stats_pcr = dpath_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = dpath_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = dpath_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = dpath_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = dpath_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = dpath_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = dpath_io_host_pcr_req_ready;
  Control ctrl(.clk(clk), .reset(reset),
       .io_dpath_sel_pc( ctrl_io_dpath_sel_pc ),
       .io_dpath_killd( ctrl_io_dpath_killd ),
       .io_dpath_ren_1( ctrl_io_dpath_ren_1 ),
       .io_dpath_ren_0( ctrl_io_dpath_ren_0 ),
       .io_dpath_sel_alu2( ctrl_io_dpath_sel_alu2 ),
       .io_dpath_sel_alu1( ctrl_io_dpath_sel_alu1 ),
       .io_dpath_sel_imm( ctrl_io_dpath_sel_imm ),
       .io_dpath_fn_dw( ctrl_io_dpath_fn_dw ),
       .io_dpath_fn_alu( ctrl_io_dpath_fn_alu ),
       .io_dpath_div_mul_val( ctrl_io_dpath_div_mul_val ),
       .io_dpath_div_mul_kill( ctrl_io_dpath_div_mul_kill ),
       //.io_dpath_div_val(  )
       //.io_dpath_div_kill(  )
       .io_dpath_csr( ctrl_io_dpath_csr ),
       .io_dpath_sret( ctrl_io_dpath_sret ),
       .io_dpath_mem_load( ctrl_io_dpath_mem_load ),
       .io_dpath_wb_load( ctrl_io_dpath_wb_load ),
       .io_dpath_ex_fp_val( ctrl_io_dpath_ex_fp_val ),
       .io_dpath_mem_fp_val( ctrl_io_dpath_mem_fp_val ),
       .io_dpath_ex_wen( ctrl_io_dpath_ex_wen ),
       .io_dpath_ex_valid( ctrl_io_dpath_ex_valid ),
       .io_dpath_mem_jalr( ctrl_io_dpath_mem_jalr ),
       .io_dpath_mem_branch( ctrl_io_dpath_mem_branch ),
       .io_dpath_mem_wen( ctrl_io_dpath_mem_wen ),
       .io_dpath_wb_wen( ctrl_io_dpath_wb_wen ),
       .io_dpath_ex_mem_type( ctrl_io_dpath_ex_mem_type ),
       .io_dpath_ex_rs2_val( ctrl_io_dpath_ex_rs2_val ),
       .io_dpath_ex_rocc_val( ctrl_io_dpath_ex_rocc_val ),
       .io_dpath_mem_rocc_val( ctrl_io_dpath_mem_rocc_val ),
       .io_dpath_bypass_1( ctrl_io_dpath_bypass_1 ),
       .io_dpath_bypass_0( ctrl_io_dpath_bypass_0 ),
       .io_dpath_bypass_src_1( ctrl_io_dpath_bypass_src_1 ),
       .io_dpath_bypass_src_0( ctrl_io_dpath_bypass_src_0 ),
       .io_dpath_ll_ready( ctrl_io_dpath_ll_ready ),
       .io_dpath_retire( ctrl_io_dpath_retire ),
       .io_dpath_exception( ctrl_io_dpath_exception ),
       .io_dpath_cause( ctrl_io_dpath_cause ),
       .io_dpath_badvaddr_wen( ctrl_io_dpath_badvaddr_wen ),
       .io_dpath_inst( dpath_io_ctrl_inst ),
       //.io_dpath_jalr_eq(  )
       .io_dpath_mem_br_taken( dpath_io_ctrl_mem_br_taken ),
       .io_dpath_mem_misprediction( dpath_io_ctrl_mem_misprediction ),
       .io_dpath_div_mul_rdy( dpath_io_ctrl_div_mul_rdy ),
       .io_dpath_ll_wen( dpath_io_ctrl_ll_wen ),
       .io_dpath_ll_waddr( dpath_io_ctrl_ll_waddr ),
       .io_dpath_ex_waddr( dpath_io_ctrl_ex_waddr ),
       .io_dpath_mem_rs1_ra( dpath_io_ctrl_mem_rs1_ra ),
       .io_dpath_mem_waddr( dpath_io_ctrl_mem_waddr ),
       .io_dpath_wb_waddr( dpath_io_ctrl_wb_waddr ),
       .io_dpath_status_ip( dpath_io_ctrl_status_ip ),
       .io_dpath_status_im( dpath_io_ctrl_status_im ),
       .io_dpath_status_zero( dpath_io_ctrl_status_zero ),
       .io_dpath_status_er( dpath_io_ctrl_status_er ),
       .io_dpath_status_vm( dpath_io_ctrl_status_vm ),
       .io_dpath_status_s64( dpath_io_ctrl_status_s64 ),
       .io_dpath_status_u64( dpath_io_ctrl_status_u64 ),
       .io_dpath_status_ef( dpath_io_ctrl_status_ef ),
       .io_dpath_status_pei( dpath_io_ctrl_status_pei ),
       .io_dpath_status_ei( dpath_io_ctrl_status_ei ),
       .io_dpath_status_ps( dpath_io_ctrl_status_ps ),
       .io_dpath_status_s( dpath_io_ctrl_status_s ),
       .io_dpath_fp_sboard_clr( dpath_io_ctrl_fp_sboard_clr ),
       .io_dpath_fp_sboard_clra( dpath_io_ctrl_fp_sboard_clra ),
       .io_dpath_csr_replay( dpath_io_ctrl_csr_replay ),
       .io_imem_req_valid( ctrl_io_imem_req_valid ),
       //.io_imem_req_bits_pc(  )
       .io_imem_resp_ready( ctrl_io_imem_resp_ready ),
       .io_imem_resp_valid( io_imem_resp_valid ),
       .io_imem_resp_bits_pc( io_imem_resp_bits_pc ),
       .io_imem_resp_bits_data( io_imem_resp_bits_data ),
       .io_imem_resp_bits_xcpt_ma( io_imem_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( io_imem_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( io_imem_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( io_imem_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_target( io_imem_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( io_imem_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_index( io_imem_btb_resp_bits_bht_index ),
       .io_imem_btb_resp_bits_bht_value( io_imem_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( ctrl_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( ctrl_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( ctrl_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_target( ctrl_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( ctrl_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_index( ctrl_io_imem_btb_update_bits_prediction_bits_bht_index ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( ctrl_io_imem_btb_update_bits_prediction_bits_bht_value ),
       //.io_imem_btb_update_bits_pc(  )
       //.io_imem_btb_update_bits_target(  )
       //.io_imem_btb_update_bits_returnAddr(  )
       .io_imem_btb_update_bits_taken( ctrl_io_imem_btb_update_bits_taken ),
       .io_imem_btb_update_bits_isJump( ctrl_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isCall( ctrl_io_imem_btb_update_bits_isCall ),
       .io_imem_btb_update_bits_isReturn( ctrl_io_imem_btb_update_bits_isReturn ),
       .io_imem_btb_update_bits_incorrectTarget( ctrl_io_imem_btb_update_bits_incorrectTarget ),
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( io_imem_ptw_req_valid ),
       .io_imem_ptw_req_bits( io_imem_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       .io_imem_invalidate( ctrl_io_imem_invalidate ),
       .io_dmem_req_ready( io_dmem_req_ready ),
       .io_dmem_req_valid( ctrl_io_dmem_req_valid ),
       .io_dmem_req_bits_kill( ctrl_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_typ( ctrl_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_phys( ctrl_io_dmem_req_bits_phys ),
       //.io_dmem_req_bits_addr(  )
       //.io_dmem_req_bits_data(  )
       //.io_dmem_req_bits_tag(  )
       .io_dmem_req_bits_cmd( ctrl_io_dmem_req_bits_cmd ),
       .io_dmem_resp_valid( io_dmem_resp_valid ),
       .io_dmem_resp_bits_nack( io_dmem_resp_bits_nack ),
       .io_dmem_resp_bits_replay( io_dmem_resp_bits_replay ),
       .io_dmem_resp_bits_typ( io_dmem_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( io_dmem_resp_bits_has_data ),
       .io_dmem_resp_bits_data( io_dmem_resp_bits_data ),
       .io_dmem_resp_bits_data_subword( io_dmem_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( io_dmem_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( io_dmem_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( io_dmem_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( io_dmem_resp_bits_store_data ),
       .io_dmem_replay_next_valid( io_dmem_replay_next_valid ),
       .io_dmem_replay_next_bits( io_dmem_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( io_dmem_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( io_dmem_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( io_dmem_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( io_dmem_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       .io_dmem_ptw_req_valid( io_dmem_ptw_req_valid ),
       .io_dmem_ptw_req_bits( io_dmem_ptw_req_bits ),
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( io_dmem_ordered ),
       //.io_dtlb_val(  )
       //.io_dtlb_kill(  )
       //.io_dtlb_rdy(  )
       //.io_dtlb_miss(  )
       //.io_xcpt_dtlb_ld(  )
       //.io_xcpt_dtlb_st(  )
       //.io_fpu_valid(  )
       //.io_fpu_fcsr_rdy(  )
       //.io_fpu_nack_mem(  )
       //.io_fpu_illegal_rm(  )
       //.io_fpu_killx(  )
       //.io_fpu_killm(  )
       //.io_fpu_dec_cmd(  )
       //.io_fpu_dec_ldst(  )
       //.io_fpu_dec_wen(  )
       //.io_fpu_dec_ren1(  )
       //.io_fpu_dec_ren2(  )
       //.io_fpu_dec_ren3(  )
       //.io_fpu_dec_swap23(  )
       //.io_fpu_dec_single(  )
       //.io_fpu_dec_fromint(  )
       //.io_fpu_dec_toint(  )
       //.io_fpu_dec_fastpipe(  )
       //.io_fpu_dec_fma(  )
       //.io_fpu_dec_round(  )
       //.io_fpu_sboard_set(  )
       //.io_fpu_sboard_clr(  )
       //.io_fpu_sboard_clra(  )
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       .io_rocc_cmd_valid( ctrl_io_rocc_cmd_valid ),
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       .io_rocc_s( ctrl_io_rocc_s ),
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_write_mask( io_rocc_imem_acquire_bits_payload_write_mask ),
       .io_rocc_imem_acquire_bits_payload_subword_addr( io_rocc_imem_acquire_bits_payload_subword_addr ),
       .io_rocc_imem_acquire_bits_payload_atomic_opcode( io_rocc_imem_acquire_bits_payload_atomic_opcode ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits ),
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       .io_rocc_exception( ctrl_io_rocc_exception )
  );
  `ifndef SYNTHESIS
    assign ctrl.io_fpu_nack_mem = {1{$random}};
    assign ctrl.io_fpu_illegal_rm = {1{$random}};
    assign ctrl.io_fpu_dec_wen = {1{$random}};
    assign ctrl.io_fpu_dec_ren1 = {1{$random}};
    assign ctrl.io_fpu_dec_ren2 = {1{$random}};
    assign ctrl.io_fpu_dec_ren3 = {1{$random}};
  `endif
  Datapath dpath(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( dpath_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( dpath_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( dpath_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( dpath_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( dpath_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( dpath_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( dpath_io_host_debug_stats_pcr ),
       .io_ctrl_sel_pc( ctrl_io_dpath_sel_pc ),
       .io_ctrl_killd( ctrl_io_dpath_killd ),
       .io_ctrl_ren_1( ctrl_io_dpath_ren_1 ),
       .io_ctrl_ren_0( ctrl_io_dpath_ren_0 ),
       .io_ctrl_sel_alu2( ctrl_io_dpath_sel_alu2 ),
       .io_ctrl_sel_alu1( ctrl_io_dpath_sel_alu1 ),
       .io_ctrl_sel_imm( ctrl_io_dpath_sel_imm ),
       .io_ctrl_fn_dw( ctrl_io_dpath_fn_dw ),
       .io_ctrl_fn_alu( ctrl_io_dpath_fn_alu ),
       .io_ctrl_div_mul_val( ctrl_io_dpath_div_mul_val ),
       .io_ctrl_div_mul_kill( ctrl_io_dpath_div_mul_kill ),
       //.io_ctrl_div_val(  )
       //.io_ctrl_div_kill(  )
       .io_ctrl_csr( ctrl_io_dpath_csr ),
       .io_ctrl_sret( ctrl_io_dpath_sret ),
       .io_ctrl_mem_load( ctrl_io_dpath_mem_load ),
       .io_ctrl_wb_load( ctrl_io_dpath_wb_load ),
       .io_ctrl_ex_fp_val( ctrl_io_dpath_ex_fp_val ),
       .io_ctrl_mem_fp_val( ctrl_io_dpath_mem_fp_val ),
       .io_ctrl_ex_wen( ctrl_io_dpath_ex_wen ),
       .io_ctrl_ex_valid( ctrl_io_dpath_ex_valid ),
       .io_ctrl_mem_jalr( ctrl_io_dpath_mem_jalr ),
       .io_ctrl_mem_branch( ctrl_io_dpath_mem_branch ),
       .io_ctrl_mem_wen( ctrl_io_dpath_mem_wen ),
       .io_ctrl_wb_wen( ctrl_io_dpath_wb_wen ),
       .io_ctrl_ex_mem_type( ctrl_io_dpath_ex_mem_type ),
       .io_ctrl_ex_rs2_val( ctrl_io_dpath_ex_rs2_val ),
       .io_ctrl_ex_rocc_val( ctrl_io_dpath_ex_rocc_val ),
       .io_ctrl_mem_rocc_val( ctrl_io_dpath_mem_rocc_val ),
       .io_ctrl_bypass_1( ctrl_io_dpath_bypass_1 ),
       .io_ctrl_bypass_0( ctrl_io_dpath_bypass_0 ),
       .io_ctrl_bypass_src_1( ctrl_io_dpath_bypass_src_1 ),
       .io_ctrl_bypass_src_0( ctrl_io_dpath_bypass_src_0 ),
       .io_ctrl_ll_ready( ctrl_io_dpath_ll_ready ),
       .io_ctrl_retire( ctrl_io_dpath_retire ),
       .io_ctrl_exception( ctrl_io_dpath_exception ),
       .io_ctrl_cause( ctrl_io_dpath_cause ),
       .io_ctrl_badvaddr_wen( ctrl_io_dpath_badvaddr_wen ),
       .io_ctrl_inst( dpath_io_ctrl_inst ),
       //.io_ctrl_jalr_eq(  )
       .io_ctrl_mem_br_taken( dpath_io_ctrl_mem_br_taken ),
       .io_ctrl_mem_misprediction( dpath_io_ctrl_mem_misprediction ),
       .io_ctrl_div_mul_rdy( dpath_io_ctrl_div_mul_rdy ),
       .io_ctrl_ll_wen( dpath_io_ctrl_ll_wen ),
       .io_ctrl_ll_waddr( dpath_io_ctrl_ll_waddr ),
       .io_ctrl_ex_waddr( dpath_io_ctrl_ex_waddr ),
       .io_ctrl_mem_rs1_ra( dpath_io_ctrl_mem_rs1_ra ),
       .io_ctrl_mem_waddr( dpath_io_ctrl_mem_waddr ),
       .io_ctrl_wb_waddr( dpath_io_ctrl_wb_waddr ),
       .io_ctrl_status_ip( dpath_io_ctrl_status_ip ),
       .io_ctrl_status_im( dpath_io_ctrl_status_im ),
       .io_ctrl_status_zero( dpath_io_ctrl_status_zero ),
       .io_ctrl_status_er( dpath_io_ctrl_status_er ),
       .io_ctrl_status_vm( dpath_io_ctrl_status_vm ),
       .io_ctrl_status_s64( dpath_io_ctrl_status_s64 ),
       .io_ctrl_status_u64( dpath_io_ctrl_status_u64 ),
       .io_ctrl_status_ef( dpath_io_ctrl_status_ef ),
       .io_ctrl_status_pei( dpath_io_ctrl_status_pei ),
       .io_ctrl_status_ei( dpath_io_ctrl_status_ei ),
       .io_ctrl_status_ps( dpath_io_ctrl_status_ps ),
       .io_ctrl_status_s( dpath_io_ctrl_status_s ),
       .io_ctrl_fp_sboard_clr( dpath_io_ctrl_fp_sboard_clr ),
       .io_ctrl_fp_sboard_clra( dpath_io_ctrl_fp_sboard_clra ),
       .io_ctrl_csr_replay( dpath_io_ctrl_csr_replay ),
       .io_dmem_req_ready( io_dmem_req_ready ),
       //.io_dmem_req_valid(  )
       //.io_dmem_req_bits_kill(  )
       //.io_dmem_req_bits_typ(  )
       //.io_dmem_req_bits_phys(  )
       .io_dmem_req_bits_addr( dpath_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_data( dpath_io_dmem_req_bits_data ),
       .io_dmem_req_bits_tag( dpath_io_dmem_req_bits_tag ),
       //.io_dmem_req_bits_cmd(  )
       .io_dmem_resp_valid( io_dmem_resp_valid ),
       .io_dmem_resp_bits_nack( io_dmem_resp_bits_nack ),
       .io_dmem_resp_bits_replay( io_dmem_resp_bits_replay ),
       .io_dmem_resp_bits_typ( io_dmem_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( io_dmem_resp_bits_has_data ),
       .io_dmem_resp_bits_data( io_dmem_resp_bits_data ),
       .io_dmem_resp_bits_data_subword( io_dmem_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( io_dmem_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( io_dmem_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( io_dmem_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( io_dmem_resp_bits_store_data ),
       .io_dmem_replay_next_valid( io_dmem_replay_next_valid ),
       .io_dmem_replay_next_bits( io_dmem_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( io_dmem_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( io_dmem_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( io_dmem_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( io_dmem_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       .io_dmem_ptw_req_valid( io_dmem_ptw_req_valid ),
       .io_dmem_ptw_req_bits( io_dmem_ptw_req_bits ),
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( io_dmem_ordered ),
       .io_ptw_ptbr( dpath_io_ptw_ptbr ),
       .io_ptw_invalidate( dpath_io_ptw_invalidate ),
       .io_ptw_sret( dpath_io_ptw_sret ),
       .io_ptw_status_ip( dpath_io_ptw_status_ip ),
       .io_ptw_status_im( dpath_io_ptw_status_im ),
       .io_ptw_status_zero( dpath_io_ptw_status_zero ),
       .io_ptw_status_er( dpath_io_ptw_status_er ),
       .io_ptw_status_vm( dpath_io_ptw_status_vm ),
       .io_ptw_status_s64( dpath_io_ptw_status_s64 ),
       .io_ptw_status_u64( dpath_io_ptw_status_u64 ),
       .io_ptw_status_ef( dpath_io_ptw_status_ef ),
       .io_ptw_status_pei( dpath_io_ptw_status_pei ),
       .io_ptw_status_ei( dpath_io_ptw_status_ei ),
       .io_ptw_status_ps( dpath_io_ptw_status_ps ),
       .io_ptw_status_s( dpath_io_ptw_status_s ),
       //.io_imem_req_valid(  )
       .io_imem_req_bits_pc( dpath_io_imem_req_bits_pc ),
       //.io_imem_resp_ready(  )
       .io_imem_resp_valid( io_imem_resp_valid ),
       .io_imem_resp_bits_pc( io_imem_resp_bits_pc ),
       .io_imem_resp_bits_data( io_imem_resp_bits_data ),
       .io_imem_resp_bits_xcpt_ma( io_imem_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( io_imem_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( io_imem_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( io_imem_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_target( io_imem_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( io_imem_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_index( io_imem_btb_resp_bits_bht_index ),
       .io_imem_btb_resp_bits_bht_value( io_imem_btb_resp_bits_bht_value ),
       //.io_imem_btb_update_valid(  )
       //.io_imem_btb_update_bits_prediction_valid(  )
       //.io_imem_btb_update_bits_prediction_bits_taken(  )
       //.io_imem_btb_update_bits_prediction_bits_target(  )
       //.io_imem_btb_update_bits_prediction_bits_entry(  )
       //.io_imem_btb_update_bits_prediction_bits_bht_index(  )
       //.io_imem_btb_update_bits_prediction_bits_bht_value(  )
       .io_imem_btb_update_bits_pc( dpath_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( dpath_io_imem_btb_update_bits_target ),
       .io_imem_btb_update_bits_returnAddr( dpath_io_imem_btb_update_bits_returnAddr ),
       //.io_imem_btb_update_bits_taken(  )
       //.io_imem_btb_update_bits_isJump(  )
       //.io_imem_btb_update_bits_isCall(  )
       //.io_imem_btb_update_bits_isReturn(  )
       //.io_imem_btb_update_bits_incorrectTarget(  )
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( io_imem_ptw_req_valid ),
       .io_imem_ptw_req_bits( io_imem_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       //.io_imem_invalidate(  )
       //.io_fpu_inst(  )
       //.io_fpu_fromint_data(  )
       //.io_fpu_fcsr_rm(  )
       //.io_fpu_fcsr_flags_valid(  )
       //.io_fpu_fcsr_flags_bits(  )
       //.io_fpu_store_data(  )
       //.io_fpu_toint_data(  )
       //.io_fpu_dmem_resp_val(  )
       //.io_fpu_dmem_resp_type(  )
       //.io_fpu_dmem_resp_tag(  )
       //.io_fpu_dmem_resp_data(  )
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       .io_rocc_cmd_bits_inst_funct( dpath_io_rocc_cmd_bits_inst_funct ),
       .io_rocc_cmd_bits_inst_rs2( dpath_io_rocc_cmd_bits_inst_rs2 ),
       .io_rocc_cmd_bits_inst_rs1( dpath_io_rocc_cmd_bits_inst_rs1 ),
       .io_rocc_cmd_bits_inst_xd( dpath_io_rocc_cmd_bits_inst_xd ),
       .io_rocc_cmd_bits_inst_xs1( dpath_io_rocc_cmd_bits_inst_xs1 ),
       .io_rocc_cmd_bits_inst_xs2( dpath_io_rocc_cmd_bits_inst_xs2 ),
       .io_rocc_cmd_bits_inst_rd( dpath_io_rocc_cmd_bits_inst_rd ),
       .io_rocc_cmd_bits_inst_opcode( dpath_io_rocc_cmd_bits_inst_opcode ),
       .io_rocc_cmd_bits_rs1( dpath_io_rocc_cmd_bits_rs1 ),
       .io_rocc_cmd_bits_rs2( dpath_io_rocc_cmd_bits_rs2 ),
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_write_mask( io_rocc_imem_acquire_bits_payload_write_mask ),
       .io_rocc_imem_acquire_bits_payload_subword_addr( io_rocc_imem_acquire_bits_payload_subword_addr ),
       .io_rocc_imem_acquire_bits_payload_atomic_opcode( io_rocc_imem_acquire_bits_payload_atomic_opcode ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
  );
  `ifndef SYNTHESIS
    assign dpath.io_fpu_fcsr_flags_valid = {1{$random}};
    assign dpath.io_fpu_fcsr_flags_bits = {1{$random}};
    assign dpath.io_fpu_store_data = {2{$random}};
    assign dpath.io_fpu_toint_data = {2{$random}};
  `endif
endmodule

module BTB(input clk, input reset,
    input [42:0] io_req,
    output io_resp_valid,
    output io_resp_bits_taken,
    output[42:0] io_resp_bits_target,
    output[2:0] io_resp_bits_entry,
    output[3:0] io_resp_bits_bht_index,
    output[1:0] io_resp_bits_bht_value,
    input  io_update_valid,
    input  io_update_bits_prediction_valid,
    input  io_update_bits_prediction_bits_taken,
    input [42:0] io_update_bits_prediction_bits_target,
    input [2:0] io_update_bits_prediction_bits_entry,
    input [3:0] io_update_bits_prediction_bits_bht_index,
    input [1:0] io_update_bits_prediction_bits_bht_value,
    input [42:0] io_update_bits_pc,
    input [42:0] io_update_bits_target,
    input [42:0] io_update_bits_returnAddr,
    input  io_update_bits_taken,
    input  io_update_bits_isJump,
    input  io_update_bits_isCall,
    input  io_update_bits_isReturn,
    input  io_update_bits_incorrectTarget,
    input  io_invalidate
);

  reg[0:0] T0 = 1'b0;
  wire T1;
  wire T2;
  wire T3;
  reg [42:0] R4;
  wire[42:0] T5;
  wire T6;
  wire T7;
  wire updateTarget;
  reg  R8;
  wire T9;
  wire updateValid;
  reg  R10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  reg  R16;
  wire T17;
  wire[1:0] T18;
  wire[1:0] T19;
  reg [1:0] T20 [15:0];
  wire[1:0] T21;
  wire[1:0] T22;
  wire T23;
  wire T24;
  reg  R25;
  wire T26;
  wire T27;
  wire T28;
  reg [1:0] R29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  reg  R37;
  wire T38;
  wire T39;
  reg [3:0] R40;
  wire[3:0] T41;
  wire[3:0] T42;
  wire[3:0] T43;
  reg [3:0] R44;
  wire[3:0] T45;
  wire[3:0] T46;
  wire[2:0] T47;
  wire[3:0] T48;
  wire[2:0] T49;
  wire[1:0] T50;
  wire T51;
  wire[1:0] T52;
  wire[1:0] T53;
  wire[3:0] T54;
  wire[3:0] T55;
  wire[7:0] hits;
  wire[7:0] T56;
  wire[7:0] T57;
  wire[3:0] T58;
  wire[1:0] T59;
  wire T60;
  wire[3:0] T61;
  wire[3:0] pageHit;
  reg [3:0] pageValid;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire[3:0] pageReplEn;
  wire[3:0] tgtPageReplEn;
  wire[3:0] tgtPageRepl;
  wire[3:0] T66;
  wire[3:0] T67;
  wire T68;
  wire[3:0] idxPageUpdateOH;
  wire[3:0] idxPageRepl;
  wire[3:0] T69;
  reg [1:0] R70;
  wire[1:0] T71;
  wire[1:0] T72;
  wire[1:0] T73;
  wire T74;
  wire doPageRepl;
  wire doTgtPageRepl;
  wire T75;
  wire T76;
  wire[3:0] T77;
  wire[3:0] T78;
  wire[3:0] idxPageReplEn;
  wire doIdxPageRepl;
  wire T79;
  wire T80;
  wire[3:0] updatePageHit;
  wire[3:0] T81;
  wire[3:0] T82;
  wire[1:0] T83;
  wire T84;
  wire[29:0] T85;
  reg [42:0] R86;
  wire[42:0] T87;
  wire[29:0] T88;
  reg [29:0] pages_0 [3:0], pages_1 [3:0], pages_2 [3:0], pages_3 [3:0];
  wire[29:0] T89;
  wire[29:0] T90;
  wire[29:0] T91;
  wire[29:0] T92;
  wire T93;
  wire[3:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire[29:0] T99;
  wire T100;
  wire T101;
  wire T102;
  wire[29:0] T103;
  wire[29:0] T104;
  wire[29:0] T105;
  wire[29:0] T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire[29:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire[29:0] T116;
  wire[1:0] T117;
  wire T118;
  wire[29:0] T119;
  wire T120;
  wire[29:0] T121;
  wire T122;
  wire T123;
  wire samePage;
  wire[29:0] T124;
  wire[29:0] T125;
  wire[3:0] T126;
  wire[2:0] T127;
  wire T128;
  wire[3:0] T129;
  wire[3:0] T130;
  wire[1:0] T131;
  wire T132;
  wire[29:0] T133;
  wire[29:0] T134;
  wire T135;
  wire[29:0] T136;
  wire[1:0] T137;
  wire T138;
  wire[29:0] T139;
  wire T140;
  wire[29:0] T141;
  wire[3:0] T142;
  wire[3:0] T143;
  wire[1:0] T144;
  reg [1:0] idxPages [7:0];
  wire[1:0] T145;
  wire[1:0] T146;
  wire T147;
  wire[1:0] T148;
  wire[1:0] T149;
  wire[1:0] T150;
  wire T151;
  wire[2:0] T152;
  reg [2:0] R153;
  wire[2:0] T154;
  wire[2:0] T155;
  wire[2:0] T156;
  wire T157;
  wire T158;
  wire T159;
  reg [2:0] R160;
  wire[2:0] T161;
  wire T162;
  wire[3:0] T163;
  wire[3:0] T164;
  wire[3:0] T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire T168;
  wire[3:0] T169;
  wire[3:0] T170;
  wire[3:0] T171;
  wire[1:0] T172;
  wire T173;
  wire[3:0] T174;
  wire[3:0] T175;
  wire[3:0] T176;
  wire[1:0] T177;
  wire[3:0] T178;
  wire[1:0] T179;
  wire T180;
  wire[3:0] T181;
  wire[3:0] T182;
  wire[3:0] T183;
  wire[1:0] T184;
  wire T185;
  wire[3:0] T186;
  wire[3:0] T187;
  wire[3:0] T188;
  wire[1:0] T189;
  wire[1:0] T190;
  wire T191;
  wire[3:0] T192;
  wire[3:0] T193;
  wire[3:0] T194;
  wire[1:0] T195;
  wire T196;
  wire[3:0] T197;
  wire[3:0] T198;
  wire[3:0] T199;
  wire[1:0] T200;
  wire[7:0] T201;
  wire[7:0] T202;
  wire[7:0] T203;
  wire[3:0] T204;
  wire[1:0] T205;
  wire T206;
  wire[12:0] T207;
  wire[12:0] T208;
  reg [12:0] idxs [7:0];
  wire[12:0] T209;
  wire[12:0] T210;
  wire T211;
  wire[12:0] T212;
  wire[1:0] T213;
  wire T214;
  wire[12:0] T215;
  wire T216;
  wire[12:0] T217;
  wire[3:0] T218;
  wire[1:0] T219;
  wire T220;
  wire[12:0] T221;
  wire T222;
  wire[12:0] T223;
  wire[1:0] T224;
  wire T225;
  wire[12:0] T226;
  wire T227;
  wire[12:0] T228;
  reg [7:0] idxValid;
  wire[7:0] T229;
  wire[7:0] T230;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[7:0] T233;
  wire[7:0] T234;
  wire[7:0] T235;
  wire[7:0] T236;
  wire[3:0] T237;
  wire[1:0] T238;
  wire T239;
  wire[3:0] T240;
  wire[3:0] T241;
  wire[3:0] T242;
  wire[3:0] T243;
  wire[1:0] T244;
  reg [1:0] tgtPages [7:0];
  wire[1:0] T245;
  wire[1:0] T246;
  wire T247;
  wire[1:0] T248;
  wire[1:0] T249;
  wire[3:0] T250;
  wire[1:0] T251;
  wire T252;
  wire T253;
  wire[3:0] T254;
  wire[3:0] T255;
  wire[3:0] T256;
  wire[3:0] T257;
  wire[1:0] T258;
  wire[1:0] T259;
  wire T260;
  wire[3:0] T261;
  wire[3:0] T262;
  wire[3:0] T263;
  wire[3:0] T264;
  wire[1:0] T265;
  wire T266;
  wire[3:0] T267;
  wire[3:0] T268;
  wire[3:0] T269;
  wire[3:0] T270;
  wire[1:0] T271;
  wire[3:0] T272;
  wire[1:0] T273;
  wire T274;
  wire[3:0] T275;
  wire[3:0] T276;
  wire[3:0] T277;
  wire[3:0] T278;
  wire[1:0] T279;
  wire T280;
  wire[3:0] T281;
  wire[3:0] T282;
  wire[3:0] T283;
  wire[3:0] T284;
  wire[1:0] T285;
  wire[1:0] T286;
  wire T287;
  wire[3:0] T288;
  wire[3:0] T289;
  wire[3:0] T290;
  wire[3:0] T291;
  wire[1:0] T292;
  wire T293;
  wire[3:0] T294;
  wire[3:0] T295;
  wire[3:0] T296;
  wire[3:0] T297;
  wire[1:0] T298;
  wire[7:0] T299;
  wire[7:0] T300;
  wire[7:0] T301;
  wire[7:0] T302;
  wire T303;
  wire T304;
  wire[7:0] T305;
  wire[7:0] T306;
  wire[3:0] T307;
  wire[1:0] T308;
  wire T309;
  wire T310;
  wire[42:0] T311;
  wire[42:0] T312;
  wire[42:0] T313;
  wire[12:0] T314;
  wire[12:0] T315;
  wire[12:0] T316;
  reg [12:0] tgts [7:0];
  wire[12:0] T317;
  wire[12:0] T318;
  wire T319;
  wire[12:0] T320;
  wire[12:0] T321;
  wire[12:0] T322;
  wire T323;
  wire[12:0] T324;
  wire[12:0] T325;
  wire[12:0] T326;
  wire T327;
  wire[12:0] T328;
  wire[12:0] T329;
  wire[12:0] T330;
  wire T331;
  wire[12:0] T332;
  wire[12:0] T333;
  wire[12:0] T334;
  wire T335;
  wire[12:0] T336;
  wire[12:0] T337;
  wire[12:0] T338;
  wire T339;
  wire[12:0] T340;
  wire[12:0] T341;
  wire[12:0] T342;
  wire T343;
  wire[12:0] T344;
  wire[12:0] T345;
  wire T346;
  wire[29:0] T347;
  wire[29:0] T348;
  wire[29:0] T349;
  wire T350;
  wire[3:0] T351;
  wire[3:0] T352;
  wire T353;
  wire[3:0] T354;
  wire[3:0] T355;
  wire T356;
  wire[3:0] T357;
  wire[3:0] T358;
  wire T359;
  wire[3:0] T360;
  wire[3:0] T361;
  wire T362;
  wire[3:0] T363;
  wire[3:0] T364;
  wire T365;
  wire[3:0] T366;
  wire[3:0] T367;
  wire T368;
  wire[3:0] T369;
  wire[3:0] T370;
  wire T371;
  wire[3:0] T372;
  wire T373;
  wire[29:0] T374;
  wire[29:0] T375;
  wire[29:0] T376;
  wire T377;
  wire[29:0] T378;
  wire[29:0] T379;
  wire[29:0] T380;
  wire T381;
  wire[29:0] T382;
  wire[29:0] T383;
  wire T384;
  wire[42:0] T385;
  reg [42:0] R386;
  wire[42:0] T387;
  wire T388;
  wire T389;
  wire[1:0] T390;
  wire T391;
  wire T392;
  reg  R393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  reg [1:0] R402;
  wire[1:0] T403;
  wire[1:0] T404;
  wire[1:0] T405;
  wire[1:0] T406;
  wire[1:0] T407;
  wire T408;
  wire T409;
  wire[1:0] T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  reg [42:0] R415;
  wire[42:0] T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  reg [0:0] useRAS [7:0];
  wire T424;
  reg  R425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  reg [0:0] isJump [7:0];
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire T494;
  wire T495;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R4 = {2{$random}};
    R8 = {1{$random}};
    R10 = {1{$random}};
    R16 = {1{$random}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      T20[initvar] = {1{$random}};
    R25 = {1{$random}};
    R29 = {1{$random}};
    R37 = {1{$random}};
    R40 = {1{$random}};
    R44 = {1{$random}};
    pageValid = {1{$random}};
    R70 = {1{$random}};
    R86 = {2{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      pages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      idxPages[initvar] = {1{$random}};
    R153 = {1{$random}};
    R160 = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      idxs[initvar] = {1{$random}};
    idxValid = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      tgtPages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      tgts[initvar] = {1{$random}};
    R386 = {2{$random}};
    R393 = {1{$random}};
    R402 = {1{$random}};
    R415 = {2{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      useRAS[initvar] = {1{$random}};
    R425 = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      isJump[initvar] = {1{$random}};
  end
`endif

  assign T1 = T2 | reset;
  assign T2 = T6 | T3;
  assign T3 = io_req == R4;
  assign T5 = io_update_valid ? io_update_bits_target : R4;
  assign T6 = T7 ^ 1'h1;
  assign T7 = T12 & updateTarget;
  assign updateTarget = updateValid & R8;
  assign T9 = io_update_valid ? io_update_bits_incorrectTarget : R8;
  assign updateValid = R8 | R10;
  assign T11 = io_update_valid ? io_update_bits_prediction_valid : R10;
  assign T12 = R16 & T13;
  assign T13 = T14 ^ 1'h1;
  assign T14 = updateValid & T15;
  assign T15 = updateTarget ^ 1'h1;
  assign T17 = reset ? 1'h0 : io_update_valid;
  assign io_resp_bits_bht_value = T18;
  assign T18 = T19;
  assign T19 = T20[T42];
  always @(posedge clk)
    if (T35)
      T20[R40] <= T22;
  assign T22 = {R25, T23};
  assign T23 = T32 | T24;
  assign T24 = T27 & R25;
  assign T26 = io_update_valid ? io_update_bits_taken : R25;
  assign T27 = T31 | T28;
  assign T28 = R29[1'h0:1'h0];
  assign T30 = io_update_valid ? io_update_bits_prediction_bits_bht_value : R29;
  assign T31 = R29[1'h1:1'h1];
  assign T32 = T34 & T33;
  assign T33 = R29[1'h0:1'h0];
  assign T34 = R29[1'h1:1'h1];
  assign T35 = T39 & T36;
  assign T36 = R37 ^ 1'h1;
  assign T38 = io_update_valid ? io_update_bits_isJump : R37;
  assign T39 = R16 & R10;
  assign T41 = io_update_valid ? io_update_bits_prediction_bits_bht_index : R40;
  assign T42 = T43;
  assign T43 = T48 ^ R44;
  assign T45 = T35 ? T46 : R44;
  assign T46 = {R25, T47};
  assign T47 = R44[2'h3:1'h1];
  assign T48 = io_req[3'h5:2'h2];
  assign io_resp_bits_bht_index = T42;
  assign io_resp_bits_entry = T49;
  assign T49 = {T310, T50};
  assign T50 = {T309, T51};
  assign T51 = T52[1'h1:1'h1];
  assign T52 = T308 | T53;
  assign T53 = T54[1'h1:1'h0];
  assign T54 = T307 | T55;
  assign T55 = hits[2'h3:1'h0];
  assign hits = T201 & T56;
  assign T56 = T57;
  assign T57 = {T178, T58};
  assign T58 = {T167, T59};
  assign T59 = {T162, T60};
  assign T60 = T61 != 4'h0;
  assign T61 = T142 & pageHit;
  assign pageHit = T129 & pageValid;
  assign T62 = reset ? 4'h0 : T63;
  assign T63 = io_invalidate ? 4'h0 : T64;
  assign T64 = T128 ? T65 : pageValid;
  assign T65 = pageValid | pageReplEn;
  assign pageReplEn = idxPageReplEn | tgtPageReplEn;
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : 4'h0;
  assign tgtPageRepl = samePage ? idxPageUpdateOH : T66;
  assign T66 = T126 | T67;
  assign T67 = {3'h0, T68};
  assign T68 = idxPageUpdateOH[2'h3:2'h3];
  assign idxPageUpdateOH = T80 ? updatePageHit : idxPageRepl;
  assign idxPageRepl = T69;
  assign T69 = 1'h1 << R70;
  assign T71 = reset ? 2'h0 : T72;
  assign T72 = T74 ? T73 : R70;
  assign T73 = R70 + 2'h1;
  assign T74 = R16 & doPageRepl;
  assign doPageRepl = doIdxPageRepl | doTgtPageRepl;
  assign doTgtPageRepl = T122 & T75;
  assign T75 = T76 ^ 1'h1;
  assign T76 = T77 != 4'h0;
  assign T77 = pageHit & T78;
  assign T78 = ~ idxPageReplEn;
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : 4'h0;
  assign doIdxPageRepl = updateTarget & T79;
  assign T79 = T80 ^ 1'h1;
  assign T80 = updatePageHit != 4'h0;
  assign updatePageHit = T81 & pageValid;
  assign T81 = T82;
  assign T82 = {T117, T83};
  assign T83 = {T115, T84};
  assign T84 = T88 == T85;
  assign T85 = R86 >> 4'hd;
  assign T87 = io_update_valid ? io_update_bits_pc : R86;
  assign T88 = pages_0[2'h0] ^ pages_1[2'h0] ^ pages_2[2'h0] ^ pages_3[2'h0];
  wire [29:0] pages_w3 = pages_0[2'h3] ^ pages_1[2'h3] ^ pages_2[2'h3];
  always @(posedge clk)
    if (T95)
      pages_3[2'h3] <= T90 ^ pages_w3;
  assign T90 = T93 ? T92 : T91;
  assign T91 = R86 >> 4'hd;
  assign T92 = io_req >> 4'hd;
  assign T93 = T94 != 4'h0;
  assign T94 = idxPageUpdateOH & 4'h5;
  assign T95 = T12 & T96;
  assign T96 = T98 & T97;
  assign T97 = pageReplEn[2'h3:2'h3];
  assign T98 = T93 ? doTgtPageRepl : doIdxPageRepl;
  wire [29:0] pages_w2 = pages_0[2'h1] ^ pages_1[2'h1] ^ pages_3[2'h1];
  always @(posedge clk)
    if (T100)
      pages_2[2'h1] <= T90 ^ pages_w2;
  assign T100 = T12 & T101;
  assign T101 = T98 & T102;
  assign T102 = pageReplEn[1'h1:1'h1];
  wire [29:0] pages_w1 = pages_0[2'h2] ^ pages_2[2'h2] ^ pages_3[2'h2];
  always @(posedge clk)
    if (T107)
      pages_1[2'h2] <= T104 ^ pages_w1;
  assign T104 = T93 ? T106 : T105;
  assign T105 = io_req >> 4'hd;
  assign T106 = R86 >> 4'hd;
  assign T107 = T12 & T108;
  assign T108 = T110 & T109;
  assign T109 = pageReplEn[2'h2:2'h2];
  assign T110 = T93 ? doIdxPageRepl : doTgtPageRepl;
  wire [29:0] pages_w0 = pages_1[2'h0] ^ pages_2[2'h0] ^ pages_3[2'h0];
  always @(posedge clk)
    if (T112)
      pages_0[2'h0] <= T104 ^ pages_w0;
  assign T112 = T12 & T113;
  assign T113 = T110 & T114;
  assign T114 = pageReplEn[1'h0:1'h0];
  assign T115 = T116 == T85;
  assign T116 = pages_0[2'h1] ^ pages_1[2'h1] ^ pages_2[2'h1] ^ pages_3[2'h1];
  assign T117 = {T120, T118};
  assign T118 = T119 == T85;
  assign T119 = pages_0[2'h2] ^ pages_1[2'h2] ^ pages_2[2'h2] ^ pages_3[2'h2];
  assign T120 = T121 == T85;
  assign T121 = pages_0[2'h3] ^ pages_1[2'h3] ^ pages_2[2'h3] ^ pages_3[2'h3];
  assign T122 = updateTarget & T123;
  assign T123 = samePage ^ 1'h1;
  assign samePage = T125 == T124;
  assign T124 = io_req >> 4'hd;
  assign T125 = R86 >> 4'hd;
  assign T126 = T127 << 1'h1;
  assign T127 = idxPageUpdateOH[2'h2:1'h0];
  assign T128 = T12 & doPageRepl;
  assign T129 = T130;
  assign T130 = {T137, T131};
  assign T131 = {T135, T132};
  assign T132 = T134 == T133;
  assign T133 = io_req >> 4'hd;
  assign T134 = pages_0[2'h0] ^ pages_1[2'h0] ^ pages_2[2'h0] ^ pages_3[2'h0];
  assign T135 = T136 == T133;
  assign T136 = pages_0[2'h1] ^ pages_1[2'h1] ^ pages_2[2'h1] ^ pages_3[2'h1];
  assign T137 = {T140, T138};
  assign T138 = T139 == T133;
  assign T139 = pages_0[2'h2] ^ pages_1[2'h2] ^ pages_2[2'h2] ^ pages_3[2'h2];
  assign T140 = T141 == T133;
  assign T141 = pages_0[2'h3] ^ pages_1[2'h3] ^ pages_2[2'h3] ^ pages_3[2'h3];
  assign T142 = T143[2'h3:1'h0];
  assign T143 = 1'h1 << T144;
  assign T144 = idxPages[3'h0];
  always @(posedge clk)
    if (T7)
      idxPages[T152] <= T146;
  assign T146 = {T151, T147};
  assign T147 = T148[1'h1:1'h1];
  assign T148 = T150 | T149;
  assign T149 = idxPageUpdateOH[1'h1:1'h0];
  assign T150 = idxPageUpdateOH[2'h3:2'h2];
  assign T151 = T150 != 2'h0;
  assign T152 = R10 ? R160 : R153;
  assign T154 = reset ? 3'h0 : T155;
  assign T155 = T157 ? T156 : R153;
  assign T156 = R153 + 3'h1;
  assign T157 = T12 & T158;
  assign T158 = T159 & updateValid;
  assign T159 = R10 ^ 1'h1;
  assign T161 = io_update_valid ? io_update_bits_prediction_bits_entry : R160;
  assign T162 = T163 != 4'h0;
  assign T163 = T164 & pageHit;
  assign T164 = T165[2'h3:1'h0];
  assign T165 = 1'h1 << T166;
  assign T166 = idxPages[3'h1];
  assign T167 = {T173, T168};
  assign T168 = T169 != 4'h0;
  assign T169 = T170 & pageHit;
  assign T170 = T171[2'h3:1'h0];
  assign T171 = 1'h1 << T172;
  assign T172 = idxPages[3'h2];
  assign T173 = T174 != 4'h0;
  assign T174 = T175 & pageHit;
  assign T175 = T176[2'h3:1'h0];
  assign T176 = 1'h1 << T177;
  assign T177 = idxPages[3'h3];
  assign T178 = {T190, T179};
  assign T179 = {T185, T180};
  assign T180 = T181 != 4'h0;
  assign T181 = T182 & pageHit;
  assign T182 = T183[2'h3:1'h0];
  assign T183 = 1'h1 << T184;
  assign T184 = idxPages[3'h4];
  assign T185 = T186 != 4'h0;
  assign T186 = T187 & pageHit;
  assign T187 = T188[2'h3:1'h0];
  assign T188 = 1'h1 << T189;
  assign T189 = idxPages[3'h5];
  assign T190 = {T196, T191};
  assign T191 = T192 != 4'h0;
  assign T192 = T193 & pageHit;
  assign T193 = T194[2'h3:1'h0];
  assign T194 = 1'h1 << T195;
  assign T195 = idxPages[3'h6];
  assign T196 = T197 != 4'h0;
  assign T197 = T198 & pageHit;
  assign T198 = T199[2'h3:1'h0];
  assign T199 = 1'h1 << T200;
  assign T200 = idxPages[3'h7];
  assign T201 = idxValid & T202;
  assign T202 = T203;
  assign T203 = {T218, T204};
  assign T204 = {T213, T205};
  assign T205 = {T211, T206};
  assign T206 = T208 == T207;
  assign T207 = io_req[4'hc:1'h0];
  assign T208 = idxs[3'h0];
  always @(posedge clk)
    if (T7)
      idxs[T152] <= T210;
  assign T210 = R86[4'hc:1'h0];
  assign T211 = T212 == T207;
  assign T212 = idxs[3'h1];
  assign T213 = {T216, T214};
  assign T214 = T215 == T207;
  assign T215 = idxs[3'h2];
  assign T216 = T217 == T207;
  assign T217 = idxs[3'h3];
  assign T218 = {T224, T219};
  assign T219 = {T222, T220};
  assign T220 = T221 == T207;
  assign T221 = idxs[3'h4];
  assign T222 = T223 == T207;
  assign T223 = idxs[3'h5];
  assign T224 = {T227, T225};
  assign T225 = T226 == T207;
  assign T226 = idxs[3'h6];
  assign T227 = T228 == T207;
  assign T228 = idxs[3'h7];
  assign T229 = reset ? 8'h0 : T230;
  assign T230 = io_invalidate ? 8'h0 : T231;
  assign T231 = T12 ? T299 : T232;
  assign T232 = T12 ? T233 : idxValid;
  assign T233 = idxValid & T234;
  assign T234 = ~ T235;
  assign T235 = T236;
  assign T236 = {T272, T237};
  assign T237 = {T259, T238};
  assign T238 = {T253, T239};
  assign T239 = T240 != 4'h0;
  assign T240 = pageReplEn & T241;
  assign T241 = T142 | T242;
  assign T242 = T243[2'h3:1'h0];
  assign T243 = 1'h1 << T244;
  assign T244 = tgtPages[3'h0];
  always @(posedge clk)
    if (T7)
      tgtPages[T152] <= T246;
  assign T246 = {T252, T247};
  assign T247 = T248[1'h1:1'h1];
  assign T248 = T251 | T249;
  assign T249 = T250[1'h1:1'h0];
  assign T250 = T76 ? pageHit : tgtPageRepl;
  assign T251 = T250[2'h3:2'h2];
  assign T252 = T251 != 2'h0;
  assign T253 = T254 != 4'h0;
  assign T254 = pageReplEn & T255;
  assign T255 = T164 | T256;
  assign T256 = T257[2'h3:1'h0];
  assign T257 = 1'h1 << T258;
  assign T258 = tgtPages[3'h1];
  assign T259 = {T266, T260};
  assign T260 = T261 != 4'h0;
  assign T261 = pageReplEn & T262;
  assign T262 = T170 | T263;
  assign T263 = T264[2'h3:1'h0];
  assign T264 = 1'h1 << T265;
  assign T265 = tgtPages[3'h2];
  assign T266 = T267 != 4'h0;
  assign T267 = pageReplEn & T268;
  assign T268 = T175 | T269;
  assign T269 = T270[2'h3:1'h0];
  assign T270 = 1'h1 << T271;
  assign T271 = tgtPages[3'h3];
  assign T272 = {T286, T273};
  assign T273 = {T280, T274};
  assign T274 = T275 != 4'h0;
  assign T275 = pageReplEn & T276;
  assign T276 = T182 | T277;
  assign T277 = T278[2'h3:1'h0];
  assign T278 = 1'h1 << T279;
  assign T279 = tgtPages[3'h4];
  assign T280 = T281 != 4'h0;
  assign T281 = pageReplEn & T282;
  assign T282 = T187 | T283;
  assign T283 = T284[2'h3:1'h0];
  assign T284 = 1'h1 << T285;
  assign T285 = tgtPages[3'h5];
  assign T286 = {T293, T287};
  assign T287 = T288 != 4'h0;
  assign T288 = pageReplEn & T289;
  assign T289 = T193 | T290;
  assign T290 = T291[2'h3:1'h0];
  assign T291 = 1'h1 << T292;
  assign T292 = tgtPages[3'h6];
  assign T293 = T294 != 4'h0;
  assign T294 = pageReplEn & T295;
  assign T295 = T198 | T296;
  assign T296 = T297[2'h3:1'h0];
  assign T297 = 1'h1 << T298;
  assign T298 = tgtPages[3'h7];
  assign T299 = T305 | T300;
  assign T300 = T302 & T301;
  assign T301 = 1'h1 << T152;
  assign T302 = T303 ? 8'hff : 8'h0;
  assign T303 = T304;
  assign T304 = updateValid;
  assign T305 = T232 & T306;
  assign T306 = ~ T301;
  assign T307 = hits[3'h7:3'h4];
  assign T308 = T54[2'h3:2'h2];
  assign T309 = T308 != 2'h0;
  assign T310 = T307 != 4'h0;
  assign io_resp_bits_target = T311;
  assign T311 = T457 ? io_update_bits_returnAddr : T312;
  assign T312 = T420 ? T385 : T313;
  assign T313 = {T347, T314};
  assign T314 = T320 | T315;
  assign T315 = T319 ? T316 : 13'h0;
  assign T316 = tgts[3'h7];
  always @(posedge clk)
    if (T7)
      tgts[T152] <= T318;
  assign T318 = io_req[4'hc:1'h0];
  assign T319 = hits[3'h7:3'h7];
  assign T320 = T324 | T321;
  assign T321 = T323 ? T322 : 13'h0;
  assign T322 = tgts[3'h6];
  assign T323 = hits[3'h6:3'h6];
  assign T324 = T328 | T325;
  assign T325 = T327 ? T326 : 13'h0;
  assign T326 = tgts[3'h5];
  assign T327 = hits[3'h5:3'h5];
  assign T328 = T332 | T329;
  assign T329 = T331 ? T330 : 13'h0;
  assign T330 = tgts[3'h4];
  assign T331 = hits[3'h4:3'h4];
  assign T332 = T336 | T333;
  assign T333 = T335 ? T334 : 13'h0;
  assign T334 = tgts[3'h3];
  assign T335 = hits[2'h3:2'h3];
  assign T336 = T340 | T337;
  assign T337 = T339 ? T338 : 13'h0;
  assign T338 = tgts[3'h2];
  assign T339 = hits[2'h2:2'h2];
  assign T340 = T344 | T341;
  assign T341 = T343 ? T342 : 13'h0;
  assign T342 = tgts[3'h1];
  assign T343 = hits[1'h1:1'h1];
  assign T344 = T346 ? T345 : 13'h0;
  assign T345 = tgts[3'h0];
  assign T346 = hits[1'h0:1'h0];
  assign T347 = T374 | T348;
  assign T348 = T350 ? T349 : 30'h0;
  assign T349 = pages_0[2'h3] ^ pages_1[2'h3] ^ pages_2[2'h3] ^ pages_3[2'h3];
  assign T350 = T351[2'h3:2'h3];
  assign T351 = T354 | T352;
  assign T352 = T353 ? T296 : 4'h0;
  assign T353 = hits[3'h7:3'h7];
  assign T354 = T357 | T355;
  assign T355 = T356 ? T290 : 4'h0;
  assign T356 = hits[3'h6:3'h6];
  assign T357 = T360 | T358;
  assign T358 = T359 ? T283 : 4'h0;
  assign T359 = hits[3'h5:3'h5];
  assign T360 = T363 | T361;
  assign T361 = T362 ? T277 : 4'h0;
  assign T362 = hits[3'h4:3'h4];
  assign T363 = T366 | T364;
  assign T364 = T365 ? T269 : 4'h0;
  assign T365 = hits[2'h3:2'h3];
  assign T366 = T369 | T367;
  assign T367 = T368 ? T263 : 4'h0;
  assign T368 = hits[2'h2:2'h2];
  assign T369 = T372 | T370;
  assign T370 = T371 ? T256 : 4'h0;
  assign T371 = hits[1'h1:1'h1];
  assign T372 = T373 ? T242 : 4'h0;
  assign T373 = hits[1'h0:1'h0];
  assign T374 = T378 | T375;
  assign T375 = T377 ? T376 : 30'h0;
  assign T376 = pages_0[2'h2] ^ pages_1[2'h2] ^ pages_2[2'h2] ^ pages_3[2'h2];
  assign T377 = T351[2'h2:2'h2];
  assign T378 = T382 | T379;
  assign T379 = T381 ? T380 : 30'h0;
  assign T380 = pages_0[2'h1] ^ pages_1[2'h1] ^ pages_2[2'h1] ^ pages_3[2'h1];
  assign T381 = T351[1'h1:1'h1];
  assign T382 = T384 ? T383 : 30'h0;
  assign T383 = pages_0[2'h0] ^ pages_1[2'h0] ^ pages_2[2'h0] ^ pages_3[2'h0];
  assign T384 = T351[1'h0:1'h0];
  assign T385 = T419 ? R415 : R386;
  assign T387 = T388 ? io_update_bits_returnAddr : R386;
  assign T388 = T397 & T389;
  assign T389 = T390[1'h0:1'h0];
  assign T390 = 1'h1 << T391;
  assign T391 = T392;
  assign T392 = R393 + 1'h1;
  assign T394 = reset ? 1'h0 : T395;
  assign T395 = T399 ? T398 : T396;
  assign T396 = T397 ? T392 : R393;
  assign T397 = io_update_valid & io_update_bits_isCall;
  assign T398 = R393 - 1'h1;
  assign T399 = T411 & T400;
  assign T400 = T401 ^ 1'h1;
  assign T401 = R402 == 2'h0;
  assign T403 = reset ? 2'h0 : T404;
  assign T404 = io_invalidate ? 2'h0 : T405;
  assign T405 = T399 ? T410 : T406;
  assign T406 = T408 ? T407 : R402;
  assign T407 = R402 + 2'h1;
  assign T408 = T397 & T409;
  assign T409 = R402 < 2'h2;
  assign T410 = R402 - 2'h1;
  assign T411 = io_update_valid & T412;
  assign T412 = T414 & T413;
  assign T413 = io_update_bits_isReturn & io_update_bits_prediction_valid;
  assign T414 = io_update_bits_isCall ^ 1'h1;
  assign T416 = T417 ? io_update_bits_returnAddr : R415;
  assign T417 = T397 & T418;
  assign T418 = T390[1'h1:1'h1];
  assign T419 = R393;
  assign T420 = T455 & T421;
  assign T421 = T428 | T422;
  assign T422 = T427 ? T423 : 1'h0;
  assign T423 = useRAS[3'h7];
  always @(posedge clk)
    if (T7)
      useRAS[T152] <= R425;
  assign T426 = io_update_valid ? io_update_bits_isReturn : R425;
  assign T427 = hits[3'h7:3'h7];
  assign T428 = T432 | T429;
  assign T429 = T431 ? T430 : 1'h0;
  assign T430 = useRAS[3'h6];
  assign T431 = hits[3'h6:3'h6];
  assign T432 = T436 | T433;
  assign T433 = T435 ? T434 : 1'h0;
  assign T434 = useRAS[3'h5];
  assign T435 = hits[3'h5:3'h5];
  assign T436 = T440 | T437;
  assign T437 = T439 ? T438 : 1'h0;
  assign T438 = useRAS[3'h4];
  assign T439 = hits[3'h4:3'h4];
  assign T440 = T444 | T441;
  assign T441 = T443 ? T442 : 1'h0;
  assign T442 = useRAS[3'h3];
  assign T443 = hits[2'h3:2'h3];
  assign T444 = T448 | T445;
  assign T445 = T447 ? T446 : 1'h0;
  assign T446 = useRAS[3'h2];
  assign T447 = hits[2'h2:2'h2];
  assign T448 = T452 | T449;
  assign T449 = T451 ? T450 : 1'h0;
  assign T450 = useRAS[3'h1];
  assign T451 = hits[1'h1:1'h1];
  assign T452 = T454 ? T453 : 1'h0;
  assign T453 = useRAS[3'h0];
  assign T454 = hits[1'h0:1'h0];
  assign T455 = T456 ^ 1'h1;
  assign T456 = R402 == 2'h0;
  assign T457 = T397 & T421;
  assign io_resp_bits_taken = T458;
  assign T458 = T459 ? 1'h0 : io_resp_valid;
  assign T459 = T493 & T460;
  assign T460 = T461 ^ 1'h1;
  assign T461 = T466 | T462;
  assign T462 = T465 ? T463 : 1'h0;
  assign T463 = isJump[3'h7];
  always @(posedge clk)
    if (T7)
      isJump[T152] <= R37;
  assign T465 = hits[3'h7:3'h7];
  assign T466 = T470 | T467;
  assign T467 = T469 ? T468 : 1'h0;
  assign T468 = isJump[3'h6];
  assign T469 = hits[3'h6:3'h6];
  assign T470 = T474 | T471;
  assign T471 = T473 ? T472 : 1'h0;
  assign T472 = isJump[3'h5];
  assign T473 = hits[3'h5:3'h5];
  assign T474 = T478 | T475;
  assign T475 = T477 ? T476 : 1'h0;
  assign T476 = isJump[3'h4];
  assign T477 = hits[3'h4:3'h4];
  assign T478 = T482 | T479;
  assign T479 = T481 ? T480 : 1'h0;
  assign T480 = isJump[3'h3];
  assign T481 = hits[2'h3:2'h3];
  assign T482 = T486 | T483;
  assign T483 = T485 ? T484 : 1'h0;
  assign T484 = isJump[3'h2];
  assign T485 = hits[2'h2:2'h2];
  assign T486 = T490 | T487;
  assign T487 = T489 ? T488 : 1'h0;
  assign T488 = isJump[3'h1];
  assign T489 = hits[1'h1:1'h1];
  assign T490 = T492 ? T491 : 1'h0;
  assign T491 = isJump[3'h0];
  assign T492 = hits[1'h0:1'h0];
  assign T493 = T494 ^ 1'h1;
  assign T494 = T18[1'h0:1'h0];
  assign io_resp_valid = T495;
  assign T495 = hits != 8'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
  if(reset) T0 <= 1'b1;
  if(!T1 && T0) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "BTB request != I$ target");
    $finish;
  end
`endif
    if(io_update_valid) begin
      R4 <= io_update_bits_target;
    end
    if(io_update_valid) begin
      R8 <= io_update_bits_incorrectTarget;
    end
    if(io_update_valid) begin
      R10 <= io_update_bits_prediction_valid;
    end
    if(reset) begin
      R16 <= 1'h0;
    end else begin
      R16 <= io_update_valid;
    end
    if(io_update_valid) begin
      R25 <= io_update_bits_taken;
    end
    if(io_update_valid) begin
      R29 <= io_update_bits_prediction_bits_bht_value;
    end
    if(io_update_valid) begin
      R37 <= io_update_bits_isJump;
    end
    if(io_update_valid) begin
      R40 <= io_update_bits_prediction_bits_bht_index;
    end
    if(T35) begin
      R44 <= T46;
    end
    if(reset) begin
      pageValid <= 4'h0;
    end else if(io_invalidate) begin
      pageValid <= 4'h0;
    end else if(T128) begin
      pageValid <= T65;
    end
    if(reset) begin
      R70 <= 2'h0;
    end else if(T74) begin
      R70 <= T73;
    end
    if(io_update_valid) begin
      R86 <= io_update_bits_pc;
    end
    if(reset) begin
      R153 <= 3'h0;
    end else if(T157) begin
      R153 <= T156;
    end
    if(io_update_valid) begin
      R160 <= io_update_bits_prediction_bits_entry;
    end
    if(reset) begin
      idxValid <= 8'h0;
    end else if(io_invalidate) begin
      idxValid <= 8'h0;
    end else if(T12) begin
      idxValid <= T299;
    end else if(T12) begin
      idxValid <= T233;
    end
    if(T388) begin
      R386 <= io_update_bits_returnAddr;
    end
    if(reset) begin
      R393 <= 1'h0;
    end else if(T399) begin
      R393 <= T398;
    end else if(T397) begin
      R393 <= T392;
    end
    if(reset) begin
      R402 <= 2'h0;
    end else if(io_invalidate) begin
      R402 <= 2'h0;
    end else if(T399) begin
      R402 <= T410;
    end else if(T408) begin
      R402 <= T407;
    end
    if(T417) begin
      R415 <= io_update_bits_returnAddr;
    end
    if(io_update_valid) begin
      R425 <= io_update_bits_isReturn;
    end
  end
endmodule

module FlowThroughSerializer_0(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [1:0] io_in_bits_header_src,
    input [1:0] io_in_bits_header_dst,
    input [511:0] io_in_bits_payload_data,
    input [3:0] io_in_bits_payload_client_xact_id,
    input [3:0] io_in_bits_payload_master_xact_id,
    input [3:0] io_in_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[3:0] io_out_bits_payload_client_xact_id,
    output[3:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[1:0] io_cnt,
    output io_done
);

  wire T0;
  wire wrap;
  reg [1:0] cnt;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg  active;
  wire T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire T12;
  wire[3:0] T13;
  reg [3:0] rbits_payload_g_type;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  reg [3:0] rbits_payload_master_xact_id;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  reg [3:0] rbits_payload_client_xact_id;
  wire[3:0] T20;
  wire[3:0] T21;
  wire[511:0] T22;
  wire[511:0] T23;
  reg [511:0] rbits_payload_data;
  wire[511:0] T24;
  wire[511:0] T25;
  wire[511:0] T26;
  wire[127:0] T27;
  wire[127:0] T28;
  wire[127:0] shifter_0;
  wire[127:0] T29;
  wire[127:0] shifter_1;
  wire[127:0] T30;
  wire T31;
  wire[1:0] T32;
  wire[127:0] T33;
  wire[127:0] shifter_2;
  wire[127:0] T34;
  wire[127:0] shifter_3;
  wire[127:0] T35;
  wire T36;
  wire T37;
  wire[1:0] T38;
  reg [1:0] rbits_header_dst;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  reg [1:0] rbits_header_src;
  wire[1:0] T42;
  wire[1:0] T43;
  wire T44;
  wire T45;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    cnt = {1{$random}};
    active = {1{$random}};
    rbits_payload_g_type = {1{$random}};
    rbits_payload_master_xact_id = {1{$random}};
    rbits_payload_client_xact_id = {1{$random}};
    rbits_payload_data = {16{$random}};
    rbits_header_dst = {1{$random}};
    rbits_header_src = {1{$random}};
  end
`endif

  assign io_done = T0;
  assign T0 = T12 & wrap;
  assign wrap = cnt == 2'h3;
  assign T1 = reset ? 2'h0 : T2;
  assign T2 = T0 ? 2'h0 : T3;
  assign T3 = T12 ? T11 : T4;
  assign T4 = T6 ? T5 : cnt;
  assign T5 = {1'h0, io_out_ready};
  assign T6 = T7 & io_in_valid;
  assign T7 = active ^ 1'h1;
  assign T8 = reset ? 1'h0 : T9;
  assign T9 = T0 ? 1'h0 : T10;
  assign T10 = T6 ? 1'h1 : active;
  assign T11 = cnt + 2'h1;
  assign T12 = active & io_out_ready;
  assign io_cnt = cnt;
  assign io_out_bits_payload_g_type = T13;
  assign T13 = active ? rbits_payload_g_type : io_in_bits_payload_g_type;
  assign T14 = reset ? io_in_bits_payload_g_type : T15;
  assign T15 = T6 ? io_in_bits_payload_g_type : rbits_payload_g_type;
  assign io_out_bits_payload_master_xact_id = T16;
  assign T16 = active ? rbits_payload_master_xact_id : io_in_bits_payload_master_xact_id;
  assign T17 = reset ? io_in_bits_payload_master_xact_id : T18;
  assign T18 = T6 ? io_in_bits_payload_master_xact_id : rbits_payload_master_xact_id;
  assign io_out_bits_payload_client_xact_id = T19;
  assign T19 = active ? rbits_payload_client_xact_id : io_in_bits_payload_client_xact_id;
  assign T20 = reset ? io_in_bits_payload_client_xact_id : T21;
  assign T21 = T6 ? io_in_bits_payload_client_xact_id : rbits_payload_client_xact_id;
  assign io_out_bits_payload_data = T22;
  assign T22 = active ? T26 : T23;
  assign T23 = active ? rbits_payload_data : io_in_bits_payload_data;
  assign T24 = reset ? io_in_bits_payload_data : T25;
  assign T25 = T6 ? io_in_bits_payload_data : rbits_payload_data;
  assign T26 = {384'h0, T27};
  assign T27 = T37 ? T33 : T28;
  assign T28 = T31 ? shifter_1 : shifter_0;
  assign shifter_0 = T29;
  assign T29 = rbits_payload_data[7'h7f:1'h0];
  assign shifter_1 = T30;
  assign T30 = rbits_payload_data[8'hff:8'h80];
  assign T31 = T32[1'h0:1'h0];
  assign T32 = cnt;
  assign T33 = T36 ? shifter_3 : shifter_2;
  assign shifter_2 = T34;
  assign T34 = rbits_payload_data[9'h17f:9'h100];
  assign shifter_3 = T35;
  assign T35 = rbits_payload_data[9'h1ff:9'h180];
  assign T36 = T32[1'h0:1'h0];
  assign T37 = T32[1'h1:1'h1];
  assign io_out_bits_header_dst = T38;
  assign T38 = active ? rbits_header_dst : io_in_bits_header_dst;
  assign T39 = reset ? io_in_bits_header_dst : T40;
  assign T40 = T6 ? io_in_bits_header_dst : rbits_header_dst;
  assign io_out_bits_header_src = T41;
  assign T41 = active ? rbits_header_src : io_in_bits_header_src;
  assign T42 = reset ? io_in_bits_header_src : T43;
  assign T43 = T6 ? io_in_bits_header_src : rbits_header_src;
  assign io_out_valid = T44;
  assign T44 = active | io_in_valid;
  assign io_in_ready = T45;
  assign T45 = active ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      cnt <= 2'h0;
    end else if(T0) begin
      cnt <= 2'h0;
    end else if(T12) begin
      cnt <= T11;
    end else if(T6) begin
      cnt <= T5;
    end
    if(reset) begin
      active <= 1'h0;
    end else if(T0) begin
      active <= 1'h0;
    end else if(T6) begin
      active <= 1'h1;
    end
    if(reset) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end else if(T6) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end
    if(reset) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end else if(T6) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end
    if(reset) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end else if(T6) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end
    if(reset) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end else if(T6) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end
    if(reset) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end else if(T6) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end
    if(reset) begin
      rbits_header_src <= io_in_bits_header_src;
    end else if(T6) begin
      rbits_header_src <= io_in_bits_header_src;
    end
  end
endmodule

module Queue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [3:0] io_enq_bits_payload_master_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[3:0] io_deq_bits_payload_master_xact_id,
    output io_count
);

  wire T0;
  wire[1:0] T1;
  reg  maybe_full;
  wire T2;
  wire T3;
  wire do_enq;
  wire T4;
  wire do_flow;
  wire T5;
  wire T6;
  wire do_deq;
  wire T7;
  wire T8;
  wire[3:0] T9;
  wire[7:0] T10;
  wire[5:0] T11;
  wire[3:0] T12;
  wire[7:0] T13;
  reg [7:0] ram [0:0];
  wire[7:0] T14;
  wire[7:0] T15;
  wire[7:0] T16;
  wire[5:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire empty;
  wire T23;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = T1[1'h0:1'h0];
  assign T1 = {maybe_full, 1'h0};
  assign T2 = reset ? 1'h0 : T3;
  assign T3 = T6 ? do_enq : maybe_full;
  assign do_enq = T5 & T4;
  assign T4 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T5 = io_enq_ready & io_enq_valid;
  assign T6 = do_enq != do_deq;
  assign do_deq = T8 & T7;
  assign T7 = do_flow ^ 1'h1;
  assign T8 = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_master_xact_id = T9;
  assign T9 = T10[2'h3:1'h0];
  assign T10 = {T19, T11};
  assign T11 = {T18, T12};
  assign T12 = T13[2'h3:1'h0];
  assign T13 = ram[1'h0];
  always @(posedge clk)
    if (do_enq)
      ram[1'h0] <= T15;
  assign T15 = T16;
  assign T16 = {io_enq_bits_header_src, T17};
  assign T17 = {io_enq_bits_header_dst, io_enq_bits_payload_master_xact_id};
  assign T18 = T13[3'h5:3'h4];
  assign T19 = T13[3'h7:3'h6];
  assign io_deq_bits_header_dst = T20;
  assign T20 = T10[3'h5:3'h4];
  assign io_deq_bits_header_src = T21;
  assign T21 = T10[3'h7:3'h6];
  assign io_deq_valid = T22;
  assign T22 = empty ^ 1'h1;
  assign empty = maybe_full ^ 1'h1;
  assign io_enq_ready = T23;
  assign T23 = maybe_full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T6) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module ICache(input clk, input reset,
    input  io_req_valid,
    input [12:0] io_req_bits_idx,
    input [18:0] io_req_bits_ppn,
    input  io_req_bits_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[31:0] io_resp_bits_data,
    output[127:0] io_resp_bits_datablock,
    input  io_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    //output[1:0] io_mem_acquire_bits_header_src
    //output[1:0] io_mem_acquire_bits_header_dst
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[3:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [3:0] io_mem_grant_bits_payload_client_xact_id,
    input [3:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[3:0] io_mem_finish_bits_payload_master_xact_id
);

  wire[3:0] FlowThroughSerializer_io_out_bits_payload_master_xact_id;
  wire[1:0] FlowThroughSerializer_io_out_bits_header_src;
  wire T0;
  wire T1;
  wire[3:0] FlowThroughSerializer_io_out_bits_payload_g_type;
  wire FlowThroughSerializer_io_done;
  wire[3:0] ack_q_io_deq_bits_payload_master_xact_id;
  wire[1:0] ack_q_io_deq_bits_header_dst;
  wire[1:0] ack_q_io_deq_bits_header_src;
  wire ack_q_io_deq_valid;
  wire FlowThroughSerializer_io_in_ready;
  wire[3:0] T2;
  wire[2:0] T3;
  wire[5:0] T4;
  wire[2:0] T5;
  wire[511:0] T6;
  wire[3:0] T7;
  wire[25:0] T8;
  wire[25:0] T9;
  reg [31:0] s2_addr;
  wire[31:0] T10;
  wire[31:0] s1_addr;
  wire[31:0] T11;
  reg [12:0] s1_pgoff;
  wire[12:0] T12;
  wire T13;
  wire rdy;
  wire T14;
  wire T15;
  wire s2_miss;
  wire T16;
  wire s2_any_tag_hit;
  wire T17;
  wire T18;
  wire s2_disparity_0;
  wire T19;
  reg  R20;
  wire T21;
  wire T22;
  wire T23;
  wire stall;
  wire T24;
  reg  s1_valid;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  reg  R31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[6:0] T37;
  wire[6:0] T38;
  wire[6:0] T39;
  wire[5:0] T40;
  wire T41;
  reg [63:0] vb_array;
  wire[63:0] T42;
  wire[127:0] T43;
  wire[127:0] T44;
  wire[127:0] T45;
  wire[127:0] T46;
  wire[127:0] T47;
  wire[127:0] T48;
  wire[127:0] T49;
  wire[127:0] T50;
  wire[6:0] T51;
  wire[5:0] T52;
  wire[127:0] T53;
  wire T54;
  wire[127:0] T55;
  wire[127:0] T56;
  wire[127:0] T57;
  wire T58;
  wire T59;
  reg  invalidated;
  wire T60;
  wire T61;
  wire T62;
  reg [1:0] state;
  wire[1:0] T63;
  wire[1:0] T64;
  wire[1:0] T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire ack_q_io_enq_ready;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire[127:0] T76;
  wire[127:0] T77;
  wire[127:0] T78;
  wire[6:0] T79;
  wire[127:0] T80;
  wire T81;
  wire[127:0] T82;
  wire[127:0] T83;
  wire[127:0] T84;
  wire T85;
  reg  s2_valid;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire s2_tag_hit_0;
  wire T92;
  reg  R93;
  wire T94;
  wire s1_tag_match_0;
  wire T95;
  wire[19:0] T96;
  wire[19:0] T97;
  wire[19:0] T98;
  wire[19:0] T99;
  reg [19:0] tag_array [63:0];
  wire[19:0] T100;
  wire[19:0] T101;
  wire[19:0] T102;
  wire[19:0] T103;
  wire[19:0] T104;
  wire[19:0] T105;
  wire[19:0] T106;
  wire[19:0] T107;
  wire[19:0] T108;
  reg [5:0] tag_raddr;
  wire[5:0] T109;
  wire[5:0] T110;
  wire[12:0] s0_pgoff;
  wire T111;
  wire T112;
  wire s0_valid;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  reg [127:0] s2_dout_0;
  wire[127:0] T121;
  wire[127:0] T122;
  reg [127:0] T123 [255:0];
  wire[127:0] T124;
  wire[127:0] T125;
  wire[511:0] FlowThroughSerializer_io_out_bits_payload_data;
  wire FlowThroughSerializer_io_out_valid;
  wire[7:0] T126;
  wire[1:0] FlowThroughSerializer_io_cnt;
  reg [7:0] R127;
  wire[7:0] T128;
  wire[7:0] T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire[31:0] T135;
  wire[127:0] T136;
  wire[6:0] T137;
  wire[1:0] T138;
  wire[5:0] T139;
  wire s2_hit;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    s2_addr = {1{$random}};
    s1_pgoff = {1{$random}};
    R20 = {1{$random}};
    s1_valid = {1{$random}};
    R31 = {1{$random}};
    vb_array = {2{$random}};
    invalidated = {1{$random}};
    state = {1{$random}};
    s2_valid = {1{$random}};
    R93 = {1{$random}};
    for (initvar = 0; initvar < 64; initvar = initvar+1)
      tag_array[initvar] = {1{$random}};
    tag_raddr = {1{$random}};
    s2_dout_0 = {4{$random}};
    for (initvar = 0; initvar < 256; initvar = initvar+1)
      T123[initvar] = {4{$random}};
    R127 = {1{$random}};
  end
`endif

  assign T0 = FlowThroughSerializer_io_done & T1;
  assign T1 = FlowThroughSerializer_io_out_bits_payload_g_type != 4'h0;
  assign io_mem_finish_bits_payload_master_xact_id = ack_q_io_deq_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = ack_q_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ack_q_io_deq_bits_header_src;
  assign io_mem_finish_valid = ack_q_io_deq_valid;
  assign io_mem_grant_ready = FlowThroughSerializer_io_in_ready;
  assign io_mem_acquire_bits_payload_atomic_opcode = T2;
  assign T2 = 4'h0;
  assign io_mem_acquire_bits_payload_subword_addr = T3;
  assign T3 = 3'h0;
  assign io_mem_acquire_bits_payload_write_mask = T4;
  assign T4 = 6'h0;
  assign io_mem_acquire_bits_payload_a_type = T5;
  assign T5 = 3'h2;
  assign io_mem_acquire_bits_payload_data = T6;
  assign T6 = 512'h0;
  assign io_mem_acquire_bits_payload_client_xact_id = T7;
  assign T7 = 4'h0;
  assign io_mem_acquire_bits_payload_addr = T8;
  assign T8 = T9;
  assign T9 = s2_addr >> 3'h6;
  assign T10 = T116 ? s1_addr : s2_addr;
  assign s1_addr = T11;
  assign T11 = {io_req_bits_ppn, s1_pgoff};
  assign T12 = T13 ? io_req_bits_idx : s1_pgoff;
  assign T13 = io_req_valid & rdy;
  assign rdy = T14;
  assign T14 = T115 & T15;
  assign T15 = s2_miss ^ 1'h1;
  assign s2_miss = s2_valid & T16;
  assign T16 = s2_any_tag_hit ^ 1'h1;
  assign s2_any_tag_hit = T17;
  assign T17 = s2_tag_hit_0 & T18;
  assign T18 = s2_disparity_0 ^ 1'h1;
  assign s2_disparity_0 = T19;
  assign T19 = R31 & R20;
  assign T21 = T22 ? 1'h0 : R20;
  assign T22 = T24 & T23;
  assign T23 = stall ^ 1'h1;
  assign stall = io_resp_ready ^ 1'h1;
  assign T24 = s1_valid & rdy;
  assign T25 = reset ? 1'h0 : T26;
  assign T26 = T30 | T27;
  assign T27 = T29 & T28;
  assign T28 = io_req_bits_kill ^ 1'h1;
  assign T29 = s1_valid & stall;
  assign T30 = io_req_valid & rdy;
  assign T32 = T22 ? T33 : R31;
  assign T33 = T34;
  assign T34 = T41 & T35;
  assign T35 = T36 - 1'h1;
  assign T36 = 1'h1 << T37;
  assign T37 = T38 + 7'h1;
  assign T38 = T39 - T39;
  assign T39 = {1'h0, T40};
  assign T40 = s1_pgoff[4'hb:3'h6];
  assign T41 = vb_array >> T39;
  assign T42 = T43[6'h3f:1'h0];
  assign T43 = reset ? 128'h0 : T44;
  assign T44 = T85 ? T76 : T45;
  assign T45 = io_invalidate ? 128'h0 : T46;
  assign T46 = T58 ? T48 : T47;
  assign T47 = {64'h0, vb_array};
  assign T48 = T55 | T49;
  assign T49 = T53 & T50;
  assign T50 = 1'h1 << T51;
  assign T51 = {1'h0, T52};
  assign T52 = s2_addr[4'hb:3'h6];
  assign T53 = T54 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T54 = 1'h1;
  assign T55 = T57 & T56;
  assign T56 = ~ T50;
  assign T57 = {64'h0, vb_array};
  assign T58 = FlowThroughSerializer_io_done & T59;
  assign T59 = invalidated ^ 1'h1;
  assign T60 = T62 ? 1'h0 : T61;
  assign T61 = io_invalidate ? 1'h1 : invalidated;
  assign T62 = 2'h0 == state;
  assign T63 = reset ? 2'h0 : T64;
  assign T64 = T74 ? 2'h0 : T65;
  assign T65 = T72 ? 2'h3 : T66;
  assign T66 = T69 ? 2'h2 : T67;
  assign T67 = T68 ? 2'h1 : state;
  assign T68 = T62 & s2_miss;
  assign T69 = T71 & T70;
  assign T70 = io_mem_acquire_ready & ack_q_io_enq_ready;
  assign T71 = 2'h1 == state;
  assign T72 = T73 & io_mem_grant_valid;
  assign T73 = 2'h2 == state;
  assign T74 = T75 & FlowThroughSerializer_io_done;
  assign T75 = 2'h3 == state;
  assign T76 = T82 | T77;
  assign T77 = T80 & T78;
  assign T78 = 1'h1 << T79;
  assign T79 = {1'h0, T52};
  assign T80 = T81 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T81 = 1'h0;
  assign T82 = T84 & T83;
  assign T83 = ~ T78;
  assign T84 = {64'h0, vb_array};
  assign T85 = s2_valid & s2_disparity_0;
  assign T86 = reset ? 1'h0 : T87;
  assign T87 = T89 | T88;
  assign T88 = io_resp_valid & stall;
  assign T89 = T91 & T90;
  assign T90 = io_req_bits_kill ^ 1'h1;
  assign T91 = s1_valid & rdy;
  assign s2_tag_hit_0 = T92;
  assign T92 = R31 & R93;
  assign T94 = T22 ? s1_tag_match_0 : R93;
  assign s1_tag_match_0 = T95;
  assign T95 = T97 == T96;
  assign T96 = s1_addr[5'h1f:4'hc];
  assign T97 = T98[5'h13:1'h0];
  assign T98 = T99[5'h13:1'h0];
  assign T99 = tag_array[tag_raddr];
  always @(posedge clk)
    if (FlowThroughSerializer_io_done)
      tag_array[T52] <= T101;
  assign T101 = T106 | T102;
  assign T102 = T105 & T103;
  assign T103 = ~ T104;
  assign T104 = 20'hfffff;
  assign T105 = tag_array[T52];
  assign T106 = T107 & T104;
  assign T107 = T108;
  assign T108 = s2_addr[5'h1f:4'hc];
  assign T109 = T112 ? T110 : tag_raddr;
  assign T110 = s0_pgoff[4'hb:3'h6];
  assign s0_pgoff = T111 ? s1_pgoff : io_req_bits_idx;
  assign T111 = s1_valid & stall;
  assign T112 = T114 & s0_valid;
  assign s0_valid = io_req_valid | T113;
  assign T113 = s1_valid & stall;
  assign T114 = FlowThroughSerializer_io_done ^ 1'h1;
  assign T115 = state == 2'h0;
  assign T116 = T118 & T117;
  assign T117 = stall ^ 1'h1;
  assign T118 = s1_valid & rdy;
  assign io_mem_acquire_valid = T119;
  assign T119 = T120 & ack_q_io_enq_ready;
  assign T120 = state == 2'h1;
  assign io_resp_bits_datablock = s2_dout_0;
  assign T121 = T132 ? T122 : s2_dout_0;
  assign T122 = T123[R127];
  always @(posedge clk)
    if (FlowThroughSerializer_io_out_valid)
      T123[T126] <= T125;
  assign T125 = FlowThroughSerializer_io_out_bits_payload_data[7'h7f:1'h0];
  assign T126 = {T52, FlowThroughSerializer_io_cnt};
  assign T128 = T130 ? T129 : R127;
  assign T129 = s0_pgoff[4'hb:3'h4];
  assign T130 = T131 & s0_valid;
  assign T131 = FlowThroughSerializer_io_out_valid ^ 1'h1;
  assign T132 = T134 & T133;
  assign T133 = stall ^ 1'h1;
  assign T134 = s1_valid & rdy;
  assign io_resp_bits_data = T135;
  assign T135 = T136[5'h1f:1'h0];
  assign T136 = s2_dout_0 >> T137;
  assign T137 = T138 << 3'h5;
  assign T138 = T139[2'h3:2'h2];
  assign T139 = s2_addr[3'h5:1'h0];
  assign io_resp_valid = s2_hit;
  assign s2_hit = s2_valid & s2_any_tag_hit;
  FlowThroughSerializer_0 FlowThroughSerializer(.clk(clk), .reset(reset),
       .io_in_ready( FlowThroughSerializer_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_header_src( io_mem_grant_bits_header_src ),
       .io_in_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_in_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_in_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_in_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_in_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_out_ready( 1'h1 ),
       .io_out_valid( FlowThroughSerializer_io_out_valid ),
       .io_out_bits_header_src( FlowThroughSerializer_io_out_bits_header_src ),
       //.io_out_bits_header_dst(  )
       .io_out_bits_payload_data( FlowThroughSerializer_io_out_bits_payload_data ),
       //.io_out_bits_payload_client_xact_id(  )
       .io_out_bits_payload_master_xact_id( FlowThroughSerializer_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( FlowThroughSerializer_io_out_bits_payload_g_type ),
       .io_cnt( FlowThroughSerializer_io_cnt ),
       .io_done( FlowThroughSerializer_io_done )
  );
  Queue_0 ack_q(.clk(clk), .reset(reset),
       .io_enq_ready( ack_q_io_enq_ready ),
       .io_enq_valid( T0 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( FlowThroughSerializer_io_out_bits_header_src ),
       .io_enq_bits_payload_master_xact_id( FlowThroughSerializer_io_out_bits_payload_master_xact_id ),
       .io_deq_ready( io_mem_finish_ready ),
       .io_deq_valid( ack_q_io_deq_valid ),
       .io_deq_bits_header_src( ack_q_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ack_q_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( ack_q_io_deq_bits_payload_master_xact_id )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign ack_q.io_enq_bits_header_src = {1{$random}};
  `endif

  always @(posedge clk) begin
    if(T116) begin
      s2_addr <= s1_addr;
    end
    if(T13) begin
      s1_pgoff <= io_req_bits_idx;
    end
    if(T22) begin
      R20 <= 1'h0;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T26;
    end
    if(T22) begin
      R31 <= T33;
    end
    vb_array <= T42;
    if(T62) begin
      invalidated <= 1'h0;
    end else if(io_invalidate) begin
      invalidated <= 1'h1;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T74) begin
      state <= 2'h0;
    end else if(T72) begin
      state <= 2'h3;
    end else if(T69) begin
      state <= 2'h2;
    end else if(T68) begin
      state <= 2'h1;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= T87;
    end
    if(T22) begin
      R93 <= s1_tag_match_0;
    end
    if(T112) begin
      tag_raddr <= T110;
    end
    if(T132) begin
      s2_dout_0 <= T122;
    end
    if(T130) begin
      R127 <= T129;
    end
  end
endmodule

module RocketCAM(input clk, input reset,
    input  io_clear,
    input  io_clear_hit,
    input [36:0] io_tag,
    output io_hit,
    output[3:0] io_hits,
    output[3:0] io_valid_bits,
    input  io_write,
    input [36:0] io_write_tag,
    input [1:0] io_write_addr
);

  reg [3:0] vb_array;
  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire T13;
  wire T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[1:0] T17;
  wire hits_0;
  wire T18;
  wire[36:0] T19;
  reg [36:0] cam_tags [3:0];
  wire[36:0] T20;
  wire T21;
  wire hits_1;
  wire T22;
  wire[36:0] T23;
  wire T24;
  wire[1:0] T25;
  wire hits_2;
  wire T26;
  wire[36:0] T27;
  wire T28;
  wire hits_3;
  wire T29;
  wire[36:0] T30;
  wire T31;
  wire T32;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    vb_array = {1{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      cam_tags[initvar] = {2{$random}};
  end
`endif

  assign io_valid_bits = vb_array;
  assign T0 = reset ? 4'h0 : T1;
  assign T1 = T13 ? T11 : T2;
  assign T2 = io_clear ? 4'h0 : T3;
  assign T3 = io_write ? T4 : vb_array;
  assign T4 = T9 | T5;
  assign T5 = T7 & T6;
  assign T6 = 1'h1 << io_write_addr;
  assign T7 = T8 ? 4'hf : 4'h0;
  assign T8 = 1'h1;
  assign T9 = vb_array & T10;
  assign T10 = ~ T6;
  assign T11 = vb_array & T12;
  assign T12 = ~ io_hits;
  assign T13 = T14 & io_clear_hit;
  assign T14 = io_clear ^ 1'h1;
  assign io_hits = T15;
  assign T15 = T16;
  assign T16 = {T25, T17};
  assign T17 = {hits_1, hits_0};
  assign hits_0 = T21 & T18;
  assign T18 = T19 == io_tag;
  assign T19 = cam_tags[2'h0];
  always @(posedge clk)
    if (io_write)
      cam_tags[io_write_addr] <= io_write_tag;
  assign T21 = vb_array[1'h0:1'h0];
  assign hits_1 = T24 & T22;
  assign T22 = T23 == io_tag;
  assign T23 = cam_tags[2'h1];
  assign T24 = vb_array[1'h1:1'h1];
  assign T25 = {hits_3, hits_2};
  assign hits_2 = T28 & T26;
  assign T26 = T27 == io_tag;
  assign T27 = cam_tags[2'h2];
  assign T28 = vb_array[2'h2:2'h2];
  assign hits_3 = T31 & T29;
  assign T29 = T30 == io_tag;
  assign T30 = cam_tags[2'h3];
  assign T31 = vb_array[2'h3:2'h3];
  assign io_hit = T32;
  assign T32 = io_hits != 4'h0;

  always @(posedge clk) begin
    if(reset) begin
      vb_array <= 4'h0;
    end else if(T13) begin
      vb_array <= T11;
    end else if(io_clear) begin
      vb_array <= 4'h0;
    end else if(io_write) begin
      vb_array <= T4;
    end
  end
endmodule

module TLB(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [6:0] io_req_bits_asid,
    input [30:0] io_req_bits_vpn,
    input  io_req_bits_passthrough,
    input  io_req_bits_instruction,
    output io_resp_miss,
    output[3:0] io_resp_hit_idx,
    output[18:0] io_resp_ppn,
    output io_resp_xcpt_ld,
    output io_resp_xcpt_st,
    output io_resp_xcpt_if,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[29:0] io_ptw_req_bits,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [18:0] io_ptw_resp_bits_ppn,
    input [5:0] io_ptw_resp_bits_perm,
    input [7:0] io_ptw_status_ip,
    input [7:0] io_ptw_status_im,
    input [6:0] io_ptw_status_zero,
    input  io_ptw_status_er,
    input  io_ptw_status_vm,
    input  io_ptw_status_s64,
    input  io_ptw_status_u64,
    input  io_ptw_status_ef,
    input  io_ptw_status_pei,
    input  io_ptw_status_ei,
    input  io_ptw_status_ps,
    input  io_ptw_status_s,
    input  io_ptw_invalidate,
    input  io_ptw_sret
);

  reg [1:0] r_refill_waddr;
  wire[1:0] T0;
  wire[1:0] repl_waddr;
  wire[1:0] T1;
  wire[2:0] T2;
  wire T3;
  wire T4;
  wire T5;
  wire[1:0] T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire T9;
  reg [3:0] R10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[6:0] T15;
  wire[1:0] T16;
  wire T17;
  wire[1:0] T18;
  wire T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire[3:0] tag_cam_io_hits;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire[3:0] T25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire[3:0] T28;
  wire[3:0] T29;
  wire T30;
  wire tlb_hit;
  wire tag_cam_io_hit;
  wire T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire T35;
  wire[3:0] T36;
  wire[3:0] tag_cam_io_valid_bits;
  wire T37;
  wire T38;
  wire has_invalid_entry;
  wire T39;
  wire T40;
  wire tlb_miss;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire[36:0] T48;
  reg [37:0] r_refill_tag;
  wire[37:0] T49;
  wire[37:0] lookup_tag;
  wire[37:0] T50;
  wire T51;
  wire T52;
  reg [1:0] state;
  wire[1:0] T53;
  wire[1:0] T54;
  wire[1:0] T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[36:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire[29:0] T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[3:0] T78;
  reg [3:0] ux_array;
  wire[3:0] T79;
  wire[3:0] T80;
  wire[3:0] T81;
  wire[3:0] T82;
  wire[3:0] T83;
  wire T84;
  wire T85;
  wire[5:0] T86;
  wire[5:0] T87;
  wire T88;
  wire T89;
  wire[3:0] T90;
  wire[3:0] T91;
  wire T92;
  wire[3:0] T93;
  reg [3:0] sx_array;
  wire[3:0] T94;
  wire[3:0] T95;
  wire[3:0] T96;
  wire[3:0] T97;
  wire[3:0] T98;
  wire T99;
  wire T100;
  wire[3:0] T101;
  wire[3:0] T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire[3:0] T108;
  reg [3:0] uw_array;
  wire[3:0] T109;
  wire[3:0] T110;
  wire[3:0] T111;
  wire[3:0] T112;
  wire[3:0] T113;
  wire T114;
  wire T115;
  wire[3:0] T116;
  wire[3:0] T117;
  wire T118;
  wire[3:0] T119;
  reg [3:0] sw_array;
  wire[3:0] T120;
  wire[3:0] T121;
  wire[3:0] T122;
  wire[3:0] T123;
  wire[3:0] T124;
  wire T125;
  wire T126;
  wire[3:0] T127;
  wire[3:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire[3:0] T134;
  reg [3:0] ur_array;
  wire[3:0] T135;
  wire[3:0] T136;
  wire[3:0] T137;
  wire[3:0] T138;
  wire[3:0] T139;
  wire T140;
  wire T141;
  wire[3:0] T142;
  wire[3:0] T143;
  wire T144;
  wire[3:0] T145;
  reg [3:0] sr_array;
  wire[3:0] T146;
  wire[3:0] T147;
  wire[3:0] T148;
  wire[3:0] T149;
  wire[3:0] T150;
  wire T151;
  wire T152;
  wire[3:0] T153;
  wire[3:0] T154;
  wire[18:0] T155;
  wire[18:0] T156;
  wire[18:0] T157;
  wire[18:0] T158;
  wire[18:0] T159;
  reg [18:0] tag_ram [3:0];
  wire[18:0] T160;
  wire T161;
  wire[18:0] T162;
  wire[18:0] T163;
  wire[18:0] T164;
  wire T165;
  wire[18:0] T166;
  wire[18:0] T167;
  wire[18:0] T168;
  wire T169;
  wire[18:0] T170;
  wire[18:0] T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    r_refill_waddr = {1{$random}};
    R10 = {1{$random}};
    r_refill_tag = {2{$random}};
    state = {1{$random}};
    ux_array = {1{$random}};
    sx_array = {1{$random}};
    uw_array = {1{$random}};
    sw_array = {1{$random}};
    ur_array = {1{$random}};
    sr_array = {1{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      tag_ram[initvar] = {1{$random}};
  end
`endif

  assign T0 = T40 ? repl_waddr : r_refill_waddr;
  assign repl_waddr = has_invalid_entry ? T32 : T1;
  assign T1 = T2[1'h1:1'h0];
  assign T2 = {T8, T3};
  assign T3 = T31 & T4;
  assign T4 = T5 - 1'h1;
  assign T5 = 1'h1 << T6;
  assign T6 = T7 + 2'h1;
  assign T7 = T8 - T8;
  assign T8 = {1'h1, T9};
  assign T9 = R10[1'h1:1'h1];
  assign T11 = T30 ? T12 : R10;
  assign T12 = T25 | T13;
  assign T13 = T24 ? 4'h0 : T14;
  assign T14 = T15[2'h3:1'h0];
  assign T15 = 4'h1 << T16;
  assign T16 = {1'h1, T17};
  assign T17 = T18[1'h1:1'h1];
  assign T18 = {T23, T19};
  assign T19 = T20[1'h1:1'h1];
  assign T20 = T22 | T21;
  assign T21 = tag_cam_io_hits[1'h1:1'h0];
  assign T22 = tag_cam_io_hits[2'h3:2'h2];
  assign T23 = T22 != 2'h0;
  assign T24 = T18[1'h0:1'h0];
  assign T25 = T27 & T26;
  assign T26 = ~ T14;
  assign T27 = T29 | T28;
  assign T28 = T17 ? 4'h0 : 4'h2;
  assign T29 = R10 & 4'hd;
  assign T30 = io_req_valid & tlb_hit;
  assign tlb_hit = io_ptw_status_vm & tag_cam_io_hit;
  assign T31 = R10 >> T8;
  assign T32 = T38 ? 1'h0 : T33;
  assign T33 = T37 ? 1'h1 : T34;
  assign T34 = T35 ? 2'h2 : 2'h3;
  assign T35 = T36[2'h2:2'h2];
  assign T36 = ~ tag_cam_io_valid_bits;
  assign T37 = T36[1'h1:1'h1];
  assign T38 = T36[1'h0:1'h0];
  assign has_invalid_entry = T39 ^ 1'h1;
  assign T39 = tag_cam_io_valid_bits == 4'hf;
  assign T40 = T47 & tlb_miss;
  assign tlb_miss = T45 & T41;
  assign T41 = T42 ^ 1'h1;
  assign T42 = T44 != T43;
  assign T43 = io_req_bits_vpn[5'h1d:5'h1d];
  assign T44 = io_req_bits_vpn[5'h1e:5'h1e];
  assign T45 = io_ptw_status_vm & T46;
  assign T46 = tag_cam_io_hit ^ 1'h1;
  assign T47 = io_req_ready & io_req_valid;
  assign T48 = r_refill_tag[6'h24:1'h0];
  assign T49 = T40 ? lookup_tag : r_refill_tag;
  assign lookup_tag = T50;
  assign T50 = {io_req_bits_asid, io_req_bits_vpn};
  assign T51 = T52 & io_ptw_resp_valid;
  assign T52 = state == 2'h2;
  assign T53 = reset ? 2'h0 : T54;
  assign T54 = io_ptw_resp_valid ? 2'h0 : T55;
  assign T55 = T64 ? 2'h3 : T56;
  assign T56 = T63 ? 2'h3 : T57;
  assign T57 = T62 ? 2'h2 : T58;
  assign T58 = T60 ? 2'h0 : T59;
  assign T59 = T40 ? 2'h1 : state;
  assign T60 = T61 & io_ptw_invalidate;
  assign T61 = state == 2'h1;
  assign T62 = T61 & io_ptw_req_ready;
  assign T63 = T62 & io_ptw_invalidate;
  assign T64 = T65 & io_ptw_invalidate;
  assign T65 = state == 2'h2;
  assign T66 = lookup_tag[6'h24:1'h0];
  assign T67 = T70 & T68;
  assign T68 = io_req_bits_instruction ? io_resp_xcpt_if : T69;
  assign T69 = io_resp_xcpt_ld & io_resp_xcpt_st;
  assign T70 = io_req_ready & io_req_valid;
  assign io_ptw_req_bits = T71;
  assign T71 = r_refill_tag[5'h1d:1'h0];
  assign io_ptw_req_valid = T72;
  assign T72 = state == 2'h1;
  assign io_resp_xcpt_if = T73;
  assign T73 = T42 | T74;
  assign T74 = tlb_hit & T75;
  assign T75 = T76 ^ 1'h1;
  assign T76 = io_ptw_status_s ? T92 : T77;
  assign T77 = T78 != 4'h0;
  assign T78 = ux_array & tag_cam_io_hits;
  assign T79 = io_ptw_resp_valid ? T80 : ux_array;
  assign T80 = T90 | T81;
  assign T81 = T83 & T82;
  assign T82 = 1'h1 << r_refill_waddr;
  assign T83 = T84 ? 4'hf : 4'h0;
  assign T84 = T85;
  assign T85 = T86[2'h2:2'h2];
  assign T86 = T87 & io_ptw_resp_bits_perm;
  assign T87 = T88 ? 6'h3f : 6'h0;
  assign T88 = T89;
  assign T89 = io_ptw_resp_bits_error ^ 1'h1;
  assign T90 = ux_array & T91;
  assign T91 = ~ T82;
  assign T92 = T93 != 4'h0;
  assign T93 = sx_array & tag_cam_io_hits;
  assign T94 = io_ptw_resp_valid ? T95 : sx_array;
  assign T95 = T101 | T96;
  assign T96 = T98 & T97;
  assign T97 = 1'h1 << r_refill_waddr;
  assign T98 = T99 ? 4'hf : 4'h0;
  assign T99 = T100;
  assign T100 = T86[3'h5:3'h5];
  assign T101 = sx_array & T102;
  assign T102 = ~ T97;
  assign io_resp_xcpt_st = T103;
  assign T103 = T42 | T104;
  assign T104 = tlb_hit & T105;
  assign T105 = T106 ^ 1'h1;
  assign T106 = io_ptw_status_s ? T118 : T107;
  assign T107 = T108 != 4'h0;
  assign T108 = uw_array & tag_cam_io_hits;
  assign T109 = io_ptw_resp_valid ? T110 : uw_array;
  assign T110 = T116 | T111;
  assign T111 = T113 & T112;
  assign T112 = 1'h1 << r_refill_waddr;
  assign T113 = T114 ? 4'hf : 4'h0;
  assign T114 = T115;
  assign T115 = T86[1'h1:1'h1];
  assign T116 = uw_array & T117;
  assign T117 = ~ T112;
  assign T118 = T119 != 4'h0;
  assign T119 = sw_array & tag_cam_io_hits;
  assign T120 = io_ptw_resp_valid ? T121 : sw_array;
  assign T121 = T127 | T122;
  assign T122 = T124 & T123;
  assign T123 = 1'h1 << r_refill_waddr;
  assign T124 = T125 ? 4'hf : 4'h0;
  assign T125 = T126;
  assign T126 = T86[3'h4:3'h4];
  assign T127 = sw_array & T128;
  assign T128 = ~ T123;
  assign io_resp_xcpt_ld = T129;
  assign T129 = T42 | T130;
  assign T130 = tlb_hit & T131;
  assign T131 = T132 ^ 1'h1;
  assign T132 = io_ptw_status_s ? T144 : T133;
  assign T133 = T134 != 4'h0;
  assign T134 = ur_array & tag_cam_io_hits;
  assign T135 = io_ptw_resp_valid ? T136 : ur_array;
  assign T136 = T142 | T137;
  assign T137 = T139 & T138;
  assign T138 = 1'h1 << r_refill_waddr;
  assign T139 = T140 ? 4'hf : 4'h0;
  assign T140 = T141;
  assign T141 = T86[1'h0:1'h0];
  assign T142 = ur_array & T143;
  assign T143 = ~ T138;
  assign T144 = T145 != 4'h0;
  assign T145 = sr_array & tag_cam_io_hits;
  assign T146 = io_ptw_resp_valid ? T147 : sr_array;
  assign T147 = T153 | T148;
  assign T148 = T150 & T149;
  assign T149 = 1'h1 << r_refill_waddr;
  assign T150 = T151 ? 4'hf : 4'h0;
  assign T151 = T152;
  assign T152 = T86[2'h3:2'h3];
  assign T153 = sr_array & T154;
  assign T154 = ~ T149;
  assign io_resp_ppn = T155;
  assign T155 = T173 ? T157 : T156;
  assign T156 = io_req_bits_vpn[5'h12:1'h0];
  assign T157 = T162 | T158;
  assign T158 = T161 ? T159 : 19'h0;
  assign T159 = tag_ram[2'h3];
  always @(posedge clk)
    if (io_ptw_resp_valid)
      tag_ram[r_refill_waddr] <= io_ptw_resp_bits_ppn;
  assign T161 = tag_cam_io_hits[2'h3:2'h3];
  assign T162 = T166 | T163;
  assign T163 = T165 ? T164 : 19'h0;
  assign T164 = tag_ram[2'h2];
  assign T165 = tag_cam_io_hits[2'h2:2'h2];
  assign T166 = T170 | T167;
  assign T167 = T169 ? T168 : 19'h0;
  assign T168 = tag_ram[2'h1];
  assign T169 = tag_cam_io_hits[1'h1:1'h1];
  assign T170 = T172 ? T171 : 19'h0;
  assign T171 = tag_ram[2'h0];
  assign T172 = tag_cam_io_hits[1'h0:1'h0];
  assign T173 = io_ptw_status_vm & T174;
  assign T174 = io_req_bits_passthrough ^ 1'h1;
  assign io_resp_hit_idx = tag_cam_io_hits;
  assign io_resp_miss = tlb_miss;
  assign io_req_ready = T175;
  assign T175 = state == 2'h0;
  RocketCAM tag_cam(.clk(clk), .reset(reset),
       .io_clear( io_ptw_invalidate ),
       .io_clear_hit( T67 ),
       .io_tag( T66 ),
       .io_hit( tag_cam_io_hit ),
       .io_hits( tag_cam_io_hits ),
       .io_valid_bits( tag_cam_io_valid_bits ),
       .io_write( T51 ),
       .io_write_tag( T48 ),
       .io_write_addr( r_refill_waddr )
  );

  always @(posedge clk) begin
    if(T40) begin
      r_refill_waddr <= repl_waddr;
    end
    if(T30) begin
      R10 <= T12;
    end
    if(T40) begin
      r_refill_tag <= lookup_tag;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if(T64) begin
      state <= 2'h3;
    end else if(T63) begin
      state <= 2'h3;
    end else if(T62) begin
      state <= 2'h2;
    end else if(T60) begin
      state <= 2'h0;
    end else if(T40) begin
      state <= 2'h1;
    end
    if(io_ptw_resp_valid) begin
      ux_array <= T80;
    end
    if(io_ptw_resp_valid) begin
      sx_array <= T95;
    end
    if(io_ptw_resp_valid) begin
      uw_array <= T110;
    end
    if(io_ptw_resp_valid) begin
      sw_array <= T121;
    end
    if(io_ptw_resp_valid) begin
      ur_array <= T136;
    end
    if(io_ptw_resp_valid) begin
      sr_array <= T147;
    end
  end
endmodule

module Frontend(input clk, input reset,
    input  io_cpu_req_valid,
    input [43:0] io_cpu_req_bits_pc,
    input  io_cpu_resp_ready,
    output io_cpu_resp_valid,
    output[43:0] io_cpu_resp_bits_pc,
    output[31:0] io_cpu_resp_bits_data,
    output io_cpu_resp_bits_xcpt_ma,
    output io_cpu_resp_bits_xcpt_if,
    output io_cpu_btb_resp_valid,
    output io_cpu_btb_resp_bits_taken,
    output[42:0] io_cpu_btb_resp_bits_target,
    output[2:0] io_cpu_btb_resp_bits_entry,
    output[3:0] io_cpu_btb_resp_bits_bht_index,
    output[1:0] io_cpu_btb_resp_bits_bht_value,
    input  io_cpu_btb_update_valid,
    input  io_cpu_btb_update_bits_prediction_valid,
    input  io_cpu_btb_update_bits_prediction_bits_taken,
    input [42:0] io_cpu_btb_update_bits_prediction_bits_target,
    input [2:0] io_cpu_btb_update_bits_prediction_bits_entry,
    input [3:0] io_cpu_btb_update_bits_prediction_bits_bht_index,
    input [1:0] io_cpu_btb_update_bits_prediction_bits_bht_value,
    input [42:0] io_cpu_btb_update_bits_pc,
    input [42:0] io_cpu_btb_update_bits_target,
    input [42:0] io_cpu_btb_update_bits_returnAddr,
    input  io_cpu_btb_update_bits_taken,
    input  io_cpu_btb_update_bits_isJump,
    input  io_cpu_btb_update_bits_isCall,
    input  io_cpu_btb_update_bits_isReturn,
    input  io_cpu_btb_update_bits_incorrectTarget,
    input  io_cpu_ptw_req_ready,
    output io_cpu_ptw_req_valid,
    output[29:0] io_cpu_ptw_req_bits,
    input  io_cpu_ptw_resp_valid,
    input  io_cpu_ptw_resp_bits_error,
    input [18:0] io_cpu_ptw_resp_bits_ppn,
    input [5:0] io_cpu_ptw_resp_bits_perm,
    input [7:0] io_cpu_ptw_status_ip,
    input [7:0] io_cpu_ptw_status_im,
    input [6:0] io_cpu_ptw_status_zero,
    input  io_cpu_ptw_status_er,
    input  io_cpu_ptw_status_vm,
    input  io_cpu_ptw_status_s64,
    input  io_cpu_ptw_status_u64,
    input  io_cpu_ptw_status_ef,
    input  io_cpu_ptw_status_pei,
    input  io_cpu_ptw_status_ei,
    input  io_cpu_ptw_status_ps,
    input  io_cpu_ptw_status_s,
    input  io_cpu_ptw_invalidate,
    input  io_cpu_ptw_sret,
    input  io_cpu_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    //output[1:0] io_mem_acquire_bits_header_src
    //output[1:0] io_mem_acquire_bits_header_dst
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[3:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [3:0] io_mem_grant_bits_payload_client_xact_id,
    input [3:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[3:0] io_mem_finish_bits_payload_master_xact_id
);

  wire[30:0] T0;
  wire[43:0] s1_pc;
  reg [43:0] s1_pc_;
  wire[43:0] T1;
  wire[43:0] T2;
  wire[43:0] npc;
  wire[43:0] T3;
  wire[43:0] predicted_npc;
  wire[43:0] pcp4;
  wire[42:0] T4;
  wire[43:0] pcp4_0;
  wire T5;
  wire T6;
  wire T7;
  wire[43:0] btbTarget;
  wire[42:0] btb_io_resp_bits_target;
  wire T8;
  wire btb_io_resp_bits_taken;
  reg [43:0] s2_pc;
  wire[43:0] T9;
  wire[43:0] T10;
  wire T11;
  wire T12;
  wire icmiss;
  wire T13;
  wire icache_io_resp_valid;
  reg  s2_valid;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire stall;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  reg  s1_same_block;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire tlb_io_resp_miss;
  wire s0_same_block;
  wire T29;
  wire[43:0] T30;
  wire[43:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire[18:0] tlb_io_resp_ppn;
  wire[12:0] T40;
  wire[43:0] T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[42:0] T46;
  wire[43:0] T47;
  wire[3:0] icache_io_mem_finish_bits_payload_master_xact_id;
  wire[1:0] icache_io_mem_finish_bits_header_dst;
  wire[1:0] icache_io_mem_finish_bits_header_src;
  wire icache_io_mem_finish_valid;
  wire icache_io_mem_grant_ready;
  wire[3:0] icache_io_mem_acquire_bits_payload_atomic_opcode;
  wire[2:0] icache_io_mem_acquire_bits_payload_subword_addr;
  wire[5:0] icache_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] icache_io_mem_acquire_bits_payload_a_type;
  wire[511:0] icache_io_mem_acquire_bits_payload_data;
  wire[3:0] icache_io_mem_acquire_bits_payload_client_xact_id;
  wire[25:0] icache_io_mem_acquire_bits_payload_addr;
  wire icache_io_mem_acquire_valid;
  wire[29:0] tlb_io_ptw_req_bits;
  wire tlb_io_ptw_req_valid;
  reg [1:0] s2_btb_resp_bits_bht_value;
  wire[1:0] T48;
  wire[1:0] btb_io_resp_bits_bht_value;
  wire T49;
  wire btb_io_resp_valid;
  reg [3:0] s2_btb_resp_bits_bht_index;
  wire[3:0] T50;
  wire[3:0] btb_io_resp_bits_bht_index;
  reg [2:0] s2_btb_resp_bits_entry;
  wire[2:0] T51;
  wire[2:0] btb_io_resp_bits_entry;
  reg [42:0] s2_btb_resp_bits_target;
  wire[42:0] T52;
  reg  s2_btb_resp_bits_taken;
  wire T53;
  reg  s2_btb_resp_valid;
  wire T54;
  wire T55;
  reg  s2_xcpt_if;
  wire T56;
  wire T57;
  wire tlb_io_resp_xcpt_if;
  wire T58;
  wire[1:0] T59;
  wire[31:0] T60;
  wire[127:0] T61;
  wire[6:0] T62;
  wire[1:0] T63;
  wire[127:0] icache_io_resp_bits_datablock;
  wire[43:0] T64;
  wire T65;
  wire T66;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    s1_pc_ = {2{$random}};
    s2_pc = {2{$random}};
    s2_valid = {1{$random}};
    s1_same_block = {1{$random}};
    s2_btb_resp_bits_bht_value = {1{$random}};
    s2_btb_resp_bits_bht_index = {1{$random}};
    s2_btb_resp_bits_entry = {1{$random}};
    s2_btb_resp_bits_target = {2{$random}};
    s2_btb_resp_bits_taken = {1{$random}};
    s2_btb_resp_valid = {1{$random}};
    s2_xcpt_if = {1{$random}};
  end
`endif

  assign T0 = s1_pc >> 4'hd;
  assign s1_pc = s1_pc_ & 44'hffffffffffe;
  assign T1 = io_cpu_req_valid ? io_cpu_req_bits_pc : T2;
  assign T2 = T18 ? npc : s1_pc_;
  assign npc = T3;
  assign T3 = icmiss ? s2_pc : predicted_npc;
  assign predicted_npc = btb_io_resp_bits_taken ? btbTarget : pcp4;
  assign pcp4 = {T5, T4};
  assign T4 = pcp4_0[6'h2a:1'h0];
  assign pcp4_0 = s1_pc + 44'h4;
  assign T5 = T7 & T6;
  assign T6 = pcp4_0[6'h2a:6'h2a];
  assign T7 = s1_pc[6'h2a:6'h2a];
  assign btbTarget = {T8, btb_io_resp_bits_target};
  assign T8 = btb_io_resp_bits_target[6'h2a:6'h2a];
  assign T9 = reset ? 44'h2000 : T10;
  assign T10 = T11 ? s1_pc : s2_pc;
  assign T11 = T18 & T12;
  assign T12 = icmiss ^ 1'h1;
  assign icmiss = s2_valid & T13;
  assign T13 = icache_io_resp_valid ^ 1'h1;
  assign T14 = reset ? 1'h1 : T15;
  assign T15 = io_cpu_req_valid ? 1'h0 : T16;
  assign T16 = T18 ? T17 : s2_valid;
  assign T17 = icmiss ^ 1'h1;
  assign T18 = stall ^ 1'h1;
  assign stall = io_cpu_resp_valid & T19;
  assign T19 = io_cpu_resp_ready ^ 1'h1;
  assign T20 = T22 & T21;
  assign T21 = icmiss ^ 1'h1;
  assign T22 = stall ^ 1'h1;
  assign T23 = T37 & T24;
  assign T24 = s1_same_block ^ 1'h1;
  assign T25 = io_cpu_req_valid ? 1'h0 : T26;
  assign T26 = T18 ? T27 : s1_same_block;
  assign T27 = s0_same_block & T28;
  assign T28 = tlb_io_resp_miss ^ 1'h1;
  assign s0_same_block = T32 & T29;
  assign T29 = T31 == T30;
  assign T30 = s1_pc & 44'h10;
  assign T31 = pcp4 & 44'h10;
  assign T32 = T34 & T33;
  assign T33 = btb_io_resp_bits_taken ^ 1'h1;
  assign T34 = T36 & T35;
  assign T35 = io_cpu_req_valid ^ 1'h1;
  assign T36 = icmiss ^ 1'h1;
  assign T37 = stall ^ 1'h1;
  assign T38 = T39 | icmiss;
  assign T39 = io_cpu_req_valid | tlb_io_resp_miss;
  assign T40 = T41[4'hc:1'h0];
  assign T41 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc;
  assign T42 = T44 & T43;
  assign T43 = s0_same_block ^ 1'h1;
  assign T44 = stall ^ 1'h1;
  assign T45 = io_cpu_invalidate | io_cpu_ptw_invalidate;
  assign T46 = T47[6'h2a:1'h0];
  assign T47 = s1_pc & 44'hffffffffffc;
  assign io_mem_finish_bits_payload_master_xact_id = icache_io_mem_finish_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = icache_io_mem_finish_bits_header_dst;
  assign io_mem_finish_bits_header_src = icache_io_mem_finish_bits_header_src;
  assign io_mem_finish_valid = icache_io_mem_finish_valid;
  assign io_mem_grant_ready = icache_io_mem_grant_ready;
  assign io_mem_acquire_bits_payload_atomic_opcode = icache_io_mem_acquire_bits_payload_atomic_opcode;
  assign io_mem_acquire_bits_payload_subword_addr = icache_io_mem_acquire_bits_payload_subword_addr;
  assign io_mem_acquire_bits_payload_write_mask = icache_io_mem_acquire_bits_payload_write_mask;
  assign io_mem_acquire_bits_payload_a_type = icache_io_mem_acquire_bits_payload_a_type;
  assign io_mem_acquire_bits_payload_data = icache_io_mem_acquire_bits_payload_data;
  assign io_mem_acquire_bits_payload_client_xact_id = icache_io_mem_acquire_bits_payload_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = icache_io_mem_acquire_bits_payload_addr;
  assign io_mem_acquire_valid = icache_io_mem_acquire_valid;
  assign io_cpu_ptw_req_bits = tlb_io_ptw_req_bits;
  assign io_cpu_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_cpu_btb_resp_bits_bht_value = s2_btb_resp_bits_bht_value;
  assign T48 = T49 ? btb_io_resp_bits_bht_value : s2_btb_resp_bits_bht_value;
  assign T49 = T11 & btb_io_resp_valid;
  assign io_cpu_btb_resp_bits_bht_index = s2_btb_resp_bits_bht_index;
  assign T50 = T49 ? btb_io_resp_bits_bht_index : s2_btb_resp_bits_bht_index;
  assign io_cpu_btb_resp_bits_entry = s2_btb_resp_bits_entry;
  assign T51 = T49 ? btb_io_resp_bits_entry : s2_btb_resp_bits_entry;
  assign io_cpu_btb_resp_bits_target = s2_btb_resp_bits_target;
  assign T52 = T49 ? btb_io_resp_bits_target : s2_btb_resp_bits_target;
  assign io_cpu_btb_resp_bits_taken = s2_btb_resp_bits_taken;
  assign T53 = T49 ? btb_io_resp_bits_taken : s2_btb_resp_bits_taken;
  assign io_cpu_btb_resp_valid = s2_btb_resp_valid;
  assign T54 = reset ? 1'h0 : T55;
  assign T55 = T11 ? btb_io_resp_valid : s2_btb_resp_valid;
  assign io_cpu_resp_bits_xcpt_if = s2_xcpt_if;
  assign T56 = reset ? 1'h0 : T57;
  assign T57 = T11 ? tlb_io_resp_xcpt_if : s2_xcpt_if;
  assign io_cpu_resp_bits_xcpt_ma = T58;
  assign T58 = T59 != 2'h0;
  assign T59 = s2_pc[1'h1:1'h0];
  assign io_cpu_resp_bits_data = T60;
  assign T60 = T61[5'h1f:1'h0];
  assign T61 = icache_io_resp_bits_datablock >> T62;
  assign T62 = T63 << 3'h5;
  assign T63 = s2_pc[2'h3:2'h2];
  assign io_cpu_resp_bits_pc = T64;
  assign T64 = s2_pc & 44'hffffffffffc;
  assign io_cpu_resp_valid = T65;
  assign T65 = s2_valid & T66;
  assign T66 = s2_xcpt_if | icache_io_resp_valid;
  BTB btb(.clk(clk), .reset(reset),
       .io_req( T46 ),
       .io_resp_valid( btb_io_resp_valid ),
       .io_resp_bits_taken( btb_io_resp_bits_taken ),
       .io_resp_bits_target( btb_io_resp_bits_target ),
       .io_resp_bits_entry( btb_io_resp_bits_entry ),
       .io_resp_bits_bht_index( btb_io_resp_bits_bht_index ),
       .io_resp_bits_bht_value( btb_io_resp_bits_bht_value ),
       .io_update_valid( io_cpu_btb_update_valid ),
       .io_update_bits_prediction_valid( io_cpu_btb_update_bits_prediction_valid ),
       .io_update_bits_prediction_bits_taken( io_cpu_btb_update_bits_prediction_bits_taken ),
       .io_update_bits_prediction_bits_target( io_cpu_btb_update_bits_prediction_bits_target ),
       .io_update_bits_prediction_bits_entry( io_cpu_btb_update_bits_prediction_bits_entry ),
       .io_update_bits_prediction_bits_bht_index( io_cpu_btb_update_bits_prediction_bits_bht_index ),
       .io_update_bits_prediction_bits_bht_value( io_cpu_btb_update_bits_prediction_bits_bht_value ),
       .io_update_bits_pc( io_cpu_btb_update_bits_pc ),
       .io_update_bits_target( io_cpu_btb_update_bits_target ),
       .io_update_bits_returnAddr( io_cpu_btb_update_bits_returnAddr ),
       .io_update_bits_taken( io_cpu_btb_update_bits_taken ),
       .io_update_bits_isJump( io_cpu_btb_update_bits_isJump ),
       .io_update_bits_isCall( io_cpu_btb_update_bits_isCall ),
       .io_update_bits_isReturn( io_cpu_btb_update_bits_isReturn ),
       .io_update_bits_incorrectTarget( io_cpu_btb_update_bits_incorrectTarget ),
       .io_invalidate( T45 )
  );
  ICache icache(.clk(clk), .reset(reset),
       .io_req_valid( T42 ),
       .io_req_bits_idx( T40 ),
       .io_req_bits_ppn( tlb_io_resp_ppn ),
       .io_req_bits_kill( T38 ),
       .io_resp_ready( T23 ),
       .io_resp_valid( icache_io_resp_valid ),
       //.io_resp_bits_data(  )
       .io_resp_bits_datablock( icache_io_resp_bits_datablock ),
       .io_invalidate( io_cpu_invalidate ),
       .io_mem_acquire_ready( io_mem_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( icache_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( icache_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( icache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( io_mem_finish_ready ),
       .io_mem_finish_valid( icache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( icache_io_mem_finish_bits_payload_master_xact_id )
  );
  TLB tlb(.clk(clk), .reset(reset),
       //.io_req_ready(  )
       .io_req_valid( T20 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T0 ),
       .io_req_bits_passthrough( 1'h0 ),
       .io_req_bits_instruction( 1'h1 ),
       .io_resp_miss( tlb_io_resp_miss ),
       //.io_resp_hit_idx(  )
       .io_resp_ppn( tlb_io_resp_ppn ),
       //.io_resp_xcpt_ld(  )
       //.io_resp_xcpt_st(  )
       .io_resp_xcpt_if( tlb_io_resp_xcpt_if ),
       .io_ptw_req_ready( io_cpu_ptw_req_ready ),
       .io_ptw_req_valid( tlb_io_ptw_req_valid ),
       .io_ptw_req_bits( tlb_io_ptw_req_bits ),
       .io_ptw_resp_valid( io_cpu_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_cpu_ptw_resp_bits_error ),
       .io_ptw_resp_bits_ppn( io_cpu_ptw_resp_bits_ppn ),
       .io_ptw_resp_bits_perm( io_cpu_ptw_resp_bits_perm ),
       .io_ptw_status_ip( io_cpu_ptw_status_ip ),
       .io_ptw_status_im( io_cpu_ptw_status_im ),
       .io_ptw_status_zero( io_cpu_ptw_status_zero ),
       .io_ptw_status_er( io_cpu_ptw_status_er ),
       .io_ptw_status_vm( io_cpu_ptw_status_vm ),
       .io_ptw_status_s64( io_cpu_ptw_status_s64 ),
       .io_ptw_status_u64( io_cpu_ptw_status_u64 ),
       .io_ptw_status_ef( io_cpu_ptw_status_ef ),
       .io_ptw_status_pei( io_cpu_ptw_status_pei ),
       .io_ptw_status_ei( io_cpu_ptw_status_ei ),
       .io_ptw_status_ps( io_cpu_ptw_status_ps ),
       .io_ptw_status_s( io_cpu_ptw_status_s ),
       .io_ptw_invalidate( io_cpu_ptw_invalidate ),
       .io_ptw_sret( io_cpu_ptw_sret )
  );

  always @(posedge clk) begin
    if(io_cpu_req_valid) begin
      s1_pc_ <= io_cpu_req_bits_pc;
    end else if(T18) begin
      s1_pc_ <= npc;
    end
    if(reset) begin
      s2_pc <= 44'h2000;
    end else if(T11) begin
      s2_pc <= s1_pc;
    end
    if(reset) begin
      s2_valid <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s2_valid <= 1'h0;
    end else if(T18) begin
      s2_valid <= T17;
    end
    if(io_cpu_req_valid) begin
      s1_same_block <= 1'h0;
    end else if(T18) begin
      s1_same_block <= T27;
    end
    if(T49) begin
      s2_btb_resp_bits_bht_value <= btb_io_resp_bits_bht_value;
    end
    if(T49) begin
      s2_btb_resp_bits_bht_index <= btb_io_resp_bits_bht_index;
    end
    if(T49) begin
      s2_btb_resp_bits_entry <= btb_io_resp_bits_entry;
    end
    if(T49) begin
      s2_btb_resp_bits_target <= btb_io_resp_bits_target;
    end
    if(T49) begin
      s2_btb_resp_bits_taken <= btb_io_resp_bits_taken;
    end
    if(reset) begin
      s2_btb_resp_valid <= 1'h0;
    end else if(T11) begin
      s2_btb_resp_valid <= btb_io_resp_valid;
    end
    if(reset) begin
      s2_xcpt_if <= 1'h0;
    end else if(T11) begin
      s2_xcpt_if <= tlb_io_resp_xcpt_if;
    end
  end
endmodule

module WritebackUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [19:0] io_req_bits_tag,
    input [5:0] io_req_bits_idx,
    input  io_req_bits_way_en,
    input [3:0] io_req_bits_client_xact_id,
    input [3:0] io_req_bits_master_xact_id,
    input [2:0] io_req_bits_r_type,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_data_req_ready,
    output io_data_req_valid,
    output io_data_req_bits_way_en,
    output[11:0] io_data_req_bits_addr,
    input [127:0] io_data_resp,
    input  io_release_ready,
    output io_release_valid,
    output[25:0] io_release_bits_addr,
    output[3:0] io_release_bits_client_xact_id,
    output[3:0] io_release_bits_master_xact_id,
    output[511:0] io_release_bits_data,
    output[2:0] io_release_bits_r_type
);

  reg [2:0] req_r_type;
  wire[2:0] T0;
  wire T1;
  reg [511:0] R2;
  wire[511:0] T3;
  wire[511:0] T4;
  wire[383:0] T5;
  wire T6;
  reg  r2_data_req_fired;
  wire T7;
  wire T8;
  reg  r1_data_req_fired;
  wire T9;
  wire T10;
  wire T11;
  reg  active;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  reg [2:0] cnt;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  reg [3:0] req_master_xact_id;
  wire[3:0] T30;
  reg [3:0] req_client_xact_id;
  wire[3:0] T31;
  wire[25:0] T32;
  wire[25:0] T33;
  reg [5:0] req_idx;
  wire[5:0] T34;
  reg [19:0] req_tag;
  wire[19:0] T35;
  wire[11:0] T36;
  wire[7:0] T37;
  wire[1:0] T38;
  reg  req_way_en;
  wire T39;
  wire fire;
  wire T40;
  wire T41;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    req_r_type = {1{$random}};
    R2 = {16{$random}};
    r2_data_req_fired = {1{$random}};
    r1_data_req_fired = {1{$random}};
    active = {1{$random}};
    cnt = {1{$random}};
    req_master_xact_id = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_idx = {1{$random}};
    req_tag = {1{$random}};
    req_way_en = {1{$random}};
  end
`endif

  assign io_release_bits_r_type = req_r_type;
  assign T0 = T1 ? io_req_bits_r_type : req_r_type;
  assign T1 = io_req_ready & io_req_valid;
  assign io_release_bits_data = R2;
  assign T3 = T6 ? T4 : R2;
  assign T4 = {io_data_resp, T5};
  assign T5 = R2[9'h1ff:8'h80];
  assign T6 = active & r2_data_req_fired;
  assign T7 = reset ? 1'h0 : T8;
  assign T8 = active ? r1_data_req_fired : r2_data_req_fired;
  assign T9 = reset ? 1'h0 : T10;
  assign T10 = T23 ? 1'h1 : T11;
  assign T11 = active ? 1'h0 : r1_data_req_fired;
  assign T12 = reset ? 1'h0 : T13;
  assign T13 = T1 ? 1'h1 : T14;
  assign T14 = T16 ? T15 : active;
  assign T15 = io_release_ready ^ 1'h1;
  assign T16 = active & T17;
  assign T17 = T27 & T18;
  assign T18 = cnt == 3'h4;
  assign T19 = reset ? 3'h0 : T20;
  assign T20 = T1 ? 3'h0 : T21;
  assign T21 = T23 ? T22 : cnt;
  assign T22 = cnt + 3'h1;
  assign T23 = active & T24;
  assign T24 = T26 & T25;
  assign T25 = io_meta_read_ready & io_meta_read_valid;
  assign T26 = io_data_req_ready & io_data_req_valid;
  assign T27 = T29 & T28;
  assign T28 = r2_data_req_fired ^ 1'h1;
  assign T29 = r1_data_req_fired ^ 1'h1;
  assign io_release_bits_master_xact_id = req_master_xact_id;
  assign T30 = T1 ? io_req_bits_master_xact_id : req_master_xact_id;
  assign io_release_bits_client_xact_id = req_client_xact_id;
  assign T31 = T1 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_release_bits_addr = T32;
  assign T32 = T33;
  assign T33 = {req_tag, req_idx};
  assign T34 = T1 ? io_req_bits_idx : req_idx;
  assign T35 = T1 ? io_req_bits_tag : req_tag;
  assign io_release_valid = T16;
  assign io_data_req_bits_addr = T36;
  assign T36 = T37 << 3'h4;
  assign T37 = {req_idx, T38};
  assign T38 = cnt[1'h1:1'h0];
  assign io_data_req_bits_way_en = req_way_en;
  assign T39 = T1 ? io_req_bits_way_en : req_way_en;
  assign io_data_req_valid = fire;
  assign fire = active & T40;
  assign T40 = cnt < 3'h4;
  assign io_meta_read_bits_tag = req_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = fire;
  assign io_req_ready = T41;
  assign T41 = active ^ 1'h1;

  always @(posedge clk) begin
    if(T1) begin
      req_r_type <= io_req_bits_r_type;
    end
    if(T6) begin
      R2 <= T4;
    end
    if(reset) begin
      r2_data_req_fired <= 1'h0;
    end else if(active) begin
      r2_data_req_fired <= r1_data_req_fired;
    end
    if(reset) begin
      r1_data_req_fired <= 1'h0;
    end else if(T23) begin
      r1_data_req_fired <= 1'h1;
    end else if(active) begin
      r1_data_req_fired <= 1'h0;
    end
    if(reset) begin
      active <= 1'h0;
    end else if(T1) begin
      active <= 1'h1;
    end else if(T16) begin
      active <= T15;
    end
    if(reset) begin
      cnt <= 3'h0;
    end else if(T1) begin
      cnt <= 3'h0;
    end else if(T23) begin
      cnt <= T22;
    end
    if(T1) begin
      req_master_xact_id <= io_req_bits_master_xact_id;
    end
    if(T1) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T1) begin
      req_idx <= io_req_bits_idx;
    end
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(T1) begin
      req_way_en <= io_req_bits_way_en;
    end
  end
endmodule

module ProbeUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [25:0] io_req_bits_addr,
    input [3:0] io_req_bits_master_xact_id,
    input [1:0] io_req_bits_p_type,
    input [3:0] io_req_bits_client_xact_id,
    input  io_rep_ready,
    output io_rep_valid,
    output[25:0] io_rep_bits_addr,
    output[3:0] io_rep_bits_client_xact_id,
    output[3:0] io_rep_bits_master_xact_id,
    output[511:0] io_rep_bits_data,
    output[2:0] io_rep_bits_r_type,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[19:0] io_wb_req_bits_tag,
    output[5:0] io_wb_req_bits_idx,
    output io_wb_req_bits_way_en,
    output[3:0] io_wb_req_bits_client_xact_id,
    output[3:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    input  io_way_en,
    input  io_mshr_rdy,
    input [1:0] io_line_state_state
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire T4;
  reg [1:0] req_p_type;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg [3:0] state;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[3:0] T28;
  wire T29;
  reg [1:0] line_state_state;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  reg  way_en;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[2:0] T43;
  wire[2:0] T44;
  wire[2:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[1:0] T50;
  wire[1:0] T51;
  wire[1:0] T52;
  reg [3:0] req_master_xact_id;
  wire[3:0] T53;
  reg [3:0] req_client_xact_id;
  wire[3:0] T54;
  wire[5:0] T55;
  reg [25:0] req_addr;
  wire[25:0] T56;
  wire[19:0] T57;
  wire T58;
  wire[1:0] T59;
  wire[1:0] T60;
  wire[1:0] T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire[19:0] T66;
  wire[5:0] T67;
  wire T68;
  wire[19:0] T69;
  wire[5:0] T70;
  wire T71;
  wire[2:0] T72;
  wire[2:0] T73;
  wire[2:0] T74;
  wire[2:0] T75;
  wire[2:0] T76;
  wire T77;
  wire T78;
  wire T79;
  wire[2:0] T80;
  wire[2:0] T81;
  wire[2:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire[1:0] T87;
  wire[1:0] T88;
  wire[1:0] T89;
  wire[511:0] T90;
  wire[3:0] T91;
  wire[3:0] T92;
  wire[25:0] T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    req_p_type = {1{$random}};
    state = {1{$random}};
    line_state_state = {1{$random}};
    way_en = {1{$random}};
    req_master_xact_id = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_addr = {1{$random}};
  end
`endif

  assign io_wb_req_bits_r_type = T0;
  assign T0 = T49 ? T43 : T1;
  assign T1 = T42 ? 3'h4 : T2;
  assign T2 = T41 ? 3'h5 : T3;
  assign T3 = T4 ? 3'h6 : 3'h4;
  assign T4 = req_p_type == 2'h2;
  assign T5 = T6 ? io_req_bits_p_type : req_p_type;
  assign T6 = T7 & io_req_valid;
  assign T7 = state == 4'h1;
  assign T8 = reset ? 4'h1 : T9;
  assign T9 = T40 ? 4'h1 : T10;
  assign T10 = T6 ? 4'h2 : T11;
  assign T11 = T38 ? 4'h3 : T12;
  assign T12 = T37 ? 4'h4 : T13;
  assign T13 = T35 ? 4'h2 : T14;
  assign T14 = T31 ? 4'h5 : T15;
  assign T15 = T32 ? T28 : T16;
  assign T16 = T26 ? 4'h1 : T17;
  assign T17 = T24 ? 4'h7 : T18;
  assign T18 = T22 ? 4'h8 : T19;
  assign T19 = T20 ? 4'h1 : state;
  assign T20 = T21 & io_meta_write_ready;
  assign T21 = state == 4'h8;
  assign T22 = T23 & io_wb_req_ready;
  assign T23 = state == 4'h7;
  assign T24 = T25 & io_wb_req_ready;
  assign T25 = state == 4'h6;
  assign T26 = T27 & io_rep_ready;
  assign T27 = state == 4'h5;
  assign T28 = T29 ? 4'h6 : 4'h8;
  assign T29 = line_state_state == 2'h3;
  assign T30 = T31 ? io_line_state_state : line_state_state;
  assign T31 = state == 4'h4;
  assign T32 = T26 & T33;
  assign T33 = way_en != 1'h0;
  assign T34 = T31 ? io_way_en : way_en;
  assign T35 = T31 & T36;
  assign T36 = io_mshr_rdy ^ 1'h1;
  assign T37 = state == 4'h3;
  assign T38 = T39 & io_meta_read_ready;
  assign T39 = state == 4'h2;
  assign T40 = state == 4'h0;
  assign T41 = req_p_type == 2'h1;
  assign T42 = req_p_type == 2'h0;
  assign T43 = T48 ? 3'h1 : T44;
  assign T44 = T47 ? 3'h2 : T45;
  assign T45 = T46 ? 3'h3 : 3'h1;
  assign T46 = req_p_type == 2'h2;
  assign T47 = req_p_type == 2'h1;
  assign T48 = req_p_type == 2'h0;
  assign T49 = T50 == 2'h3;
  assign T50 = T51[1'h1:1'h0];
  assign T51 = T33 ? line_state_state : T52;
  assign T52 = 2'h0;
  assign io_wb_req_bits_master_xact_id = req_master_xact_id;
  assign T53 = T6 ? io_req_bits_master_xact_id : req_master_xact_id;
  assign io_wb_req_bits_client_xact_id = req_client_xact_id;
  assign T54 = T6 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_wb_req_bits_way_en = way_en;
  assign io_wb_req_bits_idx = T55;
  assign T55 = req_addr[3'h5:1'h0];
  assign T56 = T6 ? io_req_bits_addr : req_addr;
  assign io_wb_req_bits_tag = T57;
  assign T57 = req_addr >> 3'h6;
  assign io_wb_req_valid = T58;
  assign T58 = state == 4'h6;
  assign io_meta_write_bits_data_coh_state = T59;
  assign T59 = T60;
  assign T60 = T65 ? 2'h0 : T61;
  assign T61 = T64 ? 2'h1 : T62;
  assign T62 = T63 ? line_state_state : line_state_state;
  assign T63 = req_p_type == 2'h2;
  assign T64 = req_p_type == 2'h1;
  assign T65 = req_p_type == 2'h0;
  assign io_meta_write_bits_data_tag = T66;
  assign T66 = req_addr >> 3'h6;
  assign io_meta_write_bits_way_en = way_en;
  assign io_meta_write_bits_idx = T67;
  assign T67 = req_addr[3'h5:1'h0];
  assign io_meta_write_valid = T68;
  assign T68 = state == 4'h8;
  assign io_meta_read_bits_tag = T69;
  assign T69 = req_addr >> 3'h6;
  assign io_meta_read_bits_idx = T70;
  assign T70 = req_addr[3'h5:1'h0];
  assign io_meta_read_valid = T71;
  assign T71 = state == 4'h2;
  assign io_rep_bits_r_type = T72;
  assign T72 = T73;
  assign T73 = T86 ? T80 : T74;
  assign T74 = T79 ? 3'h4 : T75;
  assign T75 = T78 ? 3'h5 : T76;
  assign T76 = T77 ? 3'h6 : 3'h4;
  assign T77 = req_p_type == 2'h2;
  assign T78 = req_p_type == 2'h1;
  assign T79 = req_p_type == 2'h0;
  assign T80 = T85 ? 3'h1 : T81;
  assign T81 = T84 ? 3'h2 : T82;
  assign T82 = T83 ? 3'h3 : 3'h1;
  assign T83 = req_p_type == 2'h2;
  assign T84 = req_p_type == 2'h1;
  assign T85 = req_p_type == 2'h0;
  assign T86 = T87 == 2'h3;
  assign T87 = T88[1'h1:1'h0];
  assign T88 = T33 ? line_state_state : T89;
  assign T89 = 2'h0;
  assign io_rep_bits_data = T90;
  assign T90 = 512'h0;
  assign io_rep_bits_master_xact_id = T91;
  assign T91 = req_master_xact_id;
  assign io_rep_bits_client_xact_id = T92;
  assign T92 = req_client_xact_id;
  assign io_rep_bits_addr = T93;
  assign T93 = req_addr;
  assign io_rep_valid = T94;
  assign T94 = T98 & T95;
  assign T95 = T96 ^ 1'h1;
  assign T96 = T33 & T97;
  assign T97 = line_state_state == 2'h3;
  assign T98 = state == 4'h5;
  assign io_req_ready = T99;
  assign T99 = state == 4'h1;

  always @(posedge clk) begin
    if(T6) begin
      req_p_type <= io_req_bits_p_type;
    end
    if(reset) begin
      state <= 4'h1;
    end else if(T40) begin
      state <= 4'h1;
    end else if(T6) begin
      state <= 4'h2;
    end else if(T38) begin
      state <= 4'h3;
    end else if(T37) begin
      state <= 4'h4;
    end else if(T35) begin
      state <= 4'h2;
    end else if(T31) begin
      state <= 4'h5;
    end else if(T32) begin
      state <= T28;
    end else if(T26) begin
      state <= 4'h1;
    end else if(T24) begin
      state <= 4'h7;
    end else if(T22) begin
      state <= 4'h8;
    end else if(T20) begin
      state <= 4'h1;
    end
    if(T31) begin
      line_state_state <= io_line_state_state;
    end
    if(T31) begin
      way_en <= io_way_en;
    end
    if(T6) begin
      req_master_xact_id <= io_req_bits_master_xact_id;
    end
    if(T6) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T6) begin
      req_addr <= io_req_bits_addr;
    end
  end
endmodule

module Arbiter_0(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    input [19:0] io_in_1_bits_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input [19:0] io_in_0_bits_tag,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[19:0] io_out_bits_tag,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[19:0] T2;
  wire T3;
  wire[5:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_tag = T2;
  assign T2 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign T3 = T0;
  assign io_out_bits_idx = T4;
  assign T4 = T3 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T5;
  assign T5 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T6;
  assign T6 = T7 & io_out_ready;
  assign T7 = 1'h1;
  assign io_in_1_ready = T8;
  assign T8 = T9 & io_out_ready;
  assign T9 = T10;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_1(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    input  io_in_1_bits_way_en,
    input [19:0] io_in_1_bits_data_tag,
    input [1:0] io_in_1_bits_data_coh_state,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input  io_in_0_bits_way_en,
    input [19:0] io_in_0_bits_data_tag,
    input [1:0] io_in_0_bits_data_coh_state,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output io_out_bits_way_en,
    output[19:0] io_out_bits_data_tag,
    output[1:0] io_out_bits_data_coh_state,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[1:0] T2;
  wire T3;
  wire[19:0] T4;
  wire T5;
  wire[5:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_data_coh_state = T2;
  assign T2 = T3 ? io_in_1_bits_data_coh_state : io_in_0_bits_data_coh_state;
  assign T3 = T0;
  assign io_out_bits_data_tag = T4;
  assign T4 = T3 ? io_in_1_bits_data_tag : io_in_0_bits_data_tag;
  assign io_out_bits_way_en = T5;
  assign T5 = T3 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T6;
  assign T6 = T3 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T7;
  assign T7 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T8;
  assign T8 = T9 & io_out_ready;
  assign T9 = 1'h1;
  assign io_in_1_ready = T10;
  assign T10 = T11 & io_out_ready;
  assign T11 = T12;
  assign T12 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_2(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr,
    input [3:0] io_in_1_bits_client_xact_id,
    input [511:0] io_in_1_bits_data,
    input [2:0] io_in_1_bits_a_type,
    input [5:0] io_in_1_bits_write_mask,
    input [2:0] io_in_1_bits_subword_addr,
    input [3:0] io_in_1_bits_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr,
    input [3:0] io_in_0_bits_client_xact_id,
    input [511:0] io_in_0_bits_data,
    input [2:0] io_in_0_bits_a_type,
    input [5:0] io_in_0_bits_write_mask,
    input [2:0] io_in_0_bits_subword_addr,
    input [3:0] io_in_0_bits_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr,
    output[3:0] io_out_bits_client_xact_id,
    output[511:0] io_out_bits_data,
    output[2:0] io_out_bits_a_type,
    output[5:0] io_out_bits_write_mask,
    output[2:0] io_out_bits_subword_addr,
    output[3:0] io_out_bits_atomic_opcode,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[3:0] T2;
  wire T3;
  wire[2:0] T4;
  wire[5:0] T5;
  wire[2:0] T6;
  wire[511:0] T7;
  wire[3:0] T8;
  wire[25:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_atomic_opcode = T2;
  assign T2 = T3 ? io_in_1_bits_atomic_opcode : io_in_0_bits_atomic_opcode;
  assign T3 = T0;
  assign io_out_bits_subword_addr = T4;
  assign T4 = T3 ? io_in_1_bits_subword_addr : io_in_0_bits_subword_addr;
  assign io_out_bits_write_mask = T5;
  assign T5 = T3 ? io_in_1_bits_write_mask : io_in_0_bits_write_mask;
  assign io_out_bits_a_type = T6;
  assign T6 = T3 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign io_out_bits_data = T7;
  assign T7 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_client_xact_id = T8;
  assign T8 = T3 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr = T9;
  assign T9 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T10;
  assign T10 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T11;
  assign T11 = T12 & io_out_ready;
  assign T12 = 1'h1;
  assign io_in_1_ready = T13;
  assign T13 = T14 & io_out_ready;
  assign T14 = T15;
  assign T15 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_3(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [3:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [3:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[3:0] io_out_bits_payload_master_xact_id,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[3:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_payload_master_xact_id = T2;
  assign T2 = T3 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T3 = T0;
  assign io_out_bits_header_dst = T4;
  assign T4 = T3 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T5;
  assign T5 = T3 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T6;
  assign T6 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T7;
  assign T7 = T8 & io_out_ready;
  assign T8 = 1'h1;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = T11;
  assign T11 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_4(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [19:0] io_in_1_bits_tag,
    input [5:0] io_in_1_bits_idx,
    input  io_in_1_bits_way_en,
    input [3:0] io_in_1_bits_client_xact_id,
    input [3:0] io_in_1_bits_master_xact_id,
    input [2:0] io_in_1_bits_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [19:0] io_in_0_bits_tag,
    input [5:0] io_in_0_bits_idx,
    input  io_in_0_bits_way_en,
    input [3:0] io_in_0_bits_client_xact_id,
    input [3:0] io_in_0_bits_master_xact_id,
    input [2:0] io_in_0_bits_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[19:0] io_out_bits_tag,
    output[5:0] io_out_bits_idx,
    output io_out_bits_way_en,
    output[3:0] io_out_bits_client_xact_id,
    output[3:0] io_out_bits_master_xact_id,
    output[2:0] io_out_bits_r_type,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[2:0] T2;
  wire T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire T6;
  wire[5:0] T7;
  wire[19:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_r_type = T2;
  assign T2 = T3 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign T3 = T0;
  assign io_out_bits_master_xact_id = T4;
  assign T4 = T3 ? io_in_1_bits_master_xact_id : io_in_0_bits_master_xact_id;
  assign io_out_bits_client_xact_id = T5;
  assign T5 = T3 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_way_en = T6;
  assign T6 = T3 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T7;
  assign T7 = T3 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_bits_tag = T8;
  assign T8 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_valid = T9;
  assign T9 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T10;
  assign T10 = T11 & io_out_ready;
  assign T11 = 1'h1;
  assign io_in_1_ready = T12;
  assign T12 = T13 & io_out_ready;
  assign T13 = T14;
  assign T14 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_5(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_kill,
    input [2:0] io_in_1_bits_typ,
    input  io_in_1_bits_phys,
    input [43:0] io_in_1_bits_addr,
    input [63:0] io_in_1_bits_data,
    input [7:0] io_in_1_bits_tag,
    input [4:0] io_in_1_bits_cmd,
    input [4:0] io_in_1_bits_sdq_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_kill,
    input [2:0] io_in_0_bits_typ,
    input  io_in_0_bits_phys,
    input [43:0] io_in_0_bits_addr,
    input [63:0] io_in_0_bits_data,
    input [7:0] io_in_0_bits_tag,
    input [4:0] io_in_0_bits_cmd,
    input [4:0] io_in_0_bits_sdq_id,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_kill,
    output[2:0] io_out_bits_typ,
    output io_out_bits_phys,
    output[43:0] io_out_bits_addr,
    output[63:0] io_out_bits_data,
    output[7:0] io_out_bits_tag,
    output[4:0] io_out_bits_cmd,
    output[4:0] io_out_bits_sdq_id,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[4:0] T2;
  wire T3;
  wire[4:0] T4;
  wire[7:0] T5;
  wire[63:0] T6;
  wire[43:0] T7;
  wire T8;
  wire[2:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_sdq_id = T2;
  assign T2 = T3 ? io_in_1_bits_sdq_id : io_in_0_bits_sdq_id;
  assign T3 = T0;
  assign io_out_bits_cmd = T4;
  assign T4 = T3 ? io_in_1_bits_cmd : io_in_0_bits_cmd;
  assign io_out_bits_tag = T5;
  assign T5 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_bits_data = T6;
  assign T6 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_addr = T7;
  assign T7 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_phys = T8;
  assign T8 = T3 ? io_in_1_bits_phys : io_in_0_bits_phys;
  assign io_out_bits_typ = T9;
  assign T9 = T3 ? io_in_1_bits_typ : io_in_0_bits_typ;
  assign io_out_bits_kill = T10;
  assign T10 = T3 ? io_in_1_bits_kill : io_in_0_bits_kill;
  assign io_out_valid = T11;
  assign T11 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T12;
  assign T12 = T13 & io_out_ready;
  assign T13 = 1'h1;
  assign io_in_1_ready = T14;
  assign T14 = T15 & io_out_ready;
  assign T15 = T16;
  assign T16 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_6(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits = T2;
  assign T2 = T3 ? io_in_1_bits : io_in_0_bits;
  assign T3 = T0;
  assign io_out_valid = T4;
  assign T4 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T5;
  assign T5 = T6 & io_out_ready;
  assign T6 = 1'h1;
  assign io_in_1_ready = T7;
  assign T7 = T8 & io_out_ready;
  assign T8 = T9;
  assign T9 = io_in_0_valid ^ 1'h1;
endmodule

module Queue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_kill,
    input [2:0] io_enq_bits_typ,
    input  io_enq_bits_phys,
    input [43:0] io_enq_bits_addr,
    input [63:0] io_enq_bits_data,
    input [7:0] io_enq_bits_tag,
    input [4:0] io_enq_bits_cmd,
    input [4:0] io_enq_bits_sdq_id,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_kill,
    output[2:0] io_deq_bits_typ,
    output io_deq_bits_phys,
    output[43:0] io_deq_bits_addr,
    output[63:0] io_deq_bits_data,
    output[7:0] io_deq_bits_tag,
    output[4:0] io_deq_bits_cmd,
    output[4:0] io_deq_bits_sdq_id,
    output[4:0] io_count
);

  wire[4:0] T0;
  wire[3:0] ptr_diff;
  reg [3:0] deq_ptr;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire do_deq;
  wire T4;
  wire do_flow;
  wire T5;
  reg [3:0] enq_ptr;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire do_enq;
  wire T9;
  wire T10;
  wire T11;
  wire ptr_match;
  reg  maybe_full;
  wire T12;
  wire T13;
  wire T14;
  wire[4:0] T15;
  wire[130:0] T16;
  wire[81:0] T17;
  wire[9:0] T18;
  wire[4:0] T19;
  wire[130:0] T20;
  reg [130:0] ram [15:0];
  wire[130:0] T21;
  wire[130:0] T22;
  wire[130:0] T23;
  wire[81:0] T24;
  wire[9:0] T25;
  wire[71:0] T26;
  wire[48:0] T27;
  wire[44:0] T28;
  wire[3:0] T29;
  wire[4:0] T30;
  wire[71:0] T31;
  wire[7:0] T32;
  wire[63:0] T33;
  wire[48:0] T34;
  wire[44:0] T35;
  wire[43:0] T36;
  wire T37;
  wire[3:0] T38;
  wire[2:0] T39;
  wire T40;
  wire[4:0] T41;
  wire[7:0] T42;
  wire[63:0] T43;
  wire[43:0] T44;
  wire T45;
  wire[2:0] T46;
  wire T47;
  wire T48;
  wire empty;
  wire T49;
  wire T50;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    deq_ptr = {1{$random}};
    enq_ptr = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      ram[initvar] = {5{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T11, ptr_diff};
  assign ptr_diff = enq_ptr - deq_ptr;
  assign T1 = reset ? 4'h0 : T2;
  assign T2 = do_deq ? T3 : deq_ptr;
  assign T3 = deq_ptr + 4'h1;
  assign do_deq = T5 & T4;
  assign T4 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T5 = io_deq_ready & io_deq_valid;
  assign T6 = reset ? 4'h0 : T7;
  assign T7 = do_enq ? T8 : enq_ptr;
  assign T8 = enq_ptr + 4'h1;
  assign do_enq = T10 & T9;
  assign T9 = do_flow ^ 1'h1;
  assign T10 = io_enq_ready & io_enq_valid;
  assign T11 = maybe_full & ptr_match;
  assign ptr_match = enq_ptr == deq_ptr;
  assign T12 = reset ? 1'h0 : T13;
  assign T13 = T14 ? do_enq : maybe_full;
  assign T14 = do_enq != do_deq;
  assign io_deq_bits_sdq_id = T15;
  assign T15 = T16[3'h4:1'h0];
  assign T16 = {T34, T17};
  assign T17 = {T31, T18};
  assign T18 = {T30, T19};
  assign T19 = T20[3'h4:1'h0];
  assign T20 = ram[deq_ptr];
  always @(posedge clk)
    if (do_enq)
      ram[enq_ptr] <= T22;
  assign T22 = T23;
  assign T23 = {T27, T24};
  assign T24 = {T26, T25};
  assign T25 = {io_enq_bits_cmd, io_enq_bits_sdq_id};
  assign T26 = {io_enq_bits_data, io_enq_bits_tag};
  assign T27 = {T29, T28};
  assign T28 = {io_enq_bits_phys, io_enq_bits_addr};
  assign T29 = {io_enq_bits_kill, io_enq_bits_typ};
  assign T30 = T20[4'h9:3'h5];
  assign T31 = {T33, T32};
  assign T32 = T20[5'h11:4'ha];
  assign T33 = T20[7'h51:5'h12];
  assign T34 = {T38, T35};
  assign T35 = {T37, T36};
  assign T36 = T20[7'h7d:7'h52];
  assign T37 = T20[7'h7e:7'h7e];
  assign T38 = {T40, T39};
  assign T39 = T20[8'h81:7'h7f];
  assign T40 = T20[8'h82:8'h82];
  assign io_deq_bits_cmd = T41;
  assign T41 = T16[4'h9:3'h5];
  assign io_deq_bits_tag = T42;
  assign T42 = T16[5'h11:4'ha];
  assign io_deq_bits_data = T43;
  assign T43 = T16[7'h51:5'h12];
  assign io_deq_bits_addr = T44;
  assign T44 = T16[7'h7d:7'h52];
  assign io_deq_bits_phys = T45;
  assign T45 = T16[7'h7e:7'h7e];
  assign io_deq_bits_typ = T46;
  assign T46 = T16[8'h81:7'h7f];
  assign io_deq_bits_kill = T47;
  assign T47 = T16[8'h82:8'h82];
  assign io_deq_valid = T48;
  assign T48 = empty ^ 1'h1;
  assign empty = ptr_match & T49;
  assign T49 = maybe_full ^ 1'h1;
  assign io_enq_ready = T50;
  assign T50 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      deq_ptr <= 4'h0;
    end else if(do_deq) begin
      deq_ptr <= T3;
    end
    if(reset) begin
      enq_ptr <= 4'h0;
    end else if(do_enq) begin
      enq_ptr <= T8;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T14) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module MSHR_0(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input  io_req_bits_kill,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [63:0] io_req_bits_data,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input  io_req_bits_way_en,
    input [4:0] io_req_sdq_id,
    output io_idx_match,
    output[19:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[3:0] io_mem_req_bits_client_xact_id,
    //output[511:0] io_mem_req_bits_data
    output[2:0] io_mem_req_bits_a_type,
    //output[5:0] io_mem_req_bits_write_mask
    //output[2:0] io_mem_req_bits_subword_addr
    //output[3:0] io_mem_req_bits_atomic_opcode
    output io_mem_resp_way_en,
    output[11:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[127:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[63:0] io_replay_bits_data,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [3:0] io_mem_grant_bits_payload_client_xact_id,
    input [3:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[3:0] io_mem_finish_bits_payload_master_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[19:0] io_wb_req_bits_tag,
    output[5:0] io_wb_req_bits_idx,
    output io_wb_req_bits_way_en,
    output[3:0] io_wb_req_bits_client_xact_id,
    output[3:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy
);

  wire T0;
  wire can_finish;
  wire T1;
  reg [3:0] state;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire rpq_io_deq_valid;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire refill_done;
  wire T21;
  reg [1:0] refill_count;
  wire[1:0] T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire reply;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[3:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire wb_done;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire sec_rdy;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire idx_match;
  wire[5:0] T125;
  wire[5:0] T126;
  reg [43:0] req_addr;
  wire[43:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg [1:0] meta_hazard;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  reg  req_way_en;
  wire T144;
  reg [19:0] req_old_meta_tag;
  wire[19:0] T145;
  wire T146;
  wire ackq_io_enq_ready;
  wire T147;
  wire[3:0] ackq_io_deq_bits_payload_master_xact_id;
  wire[1:0] ackq_io_deq_bits_header_dst;
  wire[1:0] ackq_io_deq_bits_header_src;
  wire T148;
  wire ackq_io_deq_valid;
  wire[4:0] rpq_io_deq_bits_sdq_id;
  wire[4:0] T149;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[7:0] rpq_io_deq_bits_tag;
  wire[63:0] rpq_io_deq_bits_data;
  wire[43:0] T150;
  wire[31:0] T151;
  wire[31:0] T152;
  wire[11:0] T153;
  wire[5:0] T154;
  wire[43:0] rpq_io_deq_bits_addr;
  wire[2:0] rpq_io_deq_bits_typ;
  wire rpq_io_deq_bits_kill;
  wire T155;
  wire T156;
  wire[1:0] T157;
  wire[1:0] T158;
  reg [1:0] line_state_state;
  wire[1:0] T159;
  wire[1:0] T160;
  wire[1:0] T161;
  wire[1:0] meta_on_grant_state;
  wire[1:0] T162;
  wire[1:0] T163;
  wire[1:0] T164;
  wire T165;
  wire[1:0] T166;
  wire T167;
  wire T168;
  wire T169;
  wire[1:0] meta_on_flush_state;
  wire[1:0] meta_on_hit_state;
  wire[1:0] T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire[127:0] T183;
  reg [63:0] req_data;
  wire[63:0] T184;
  wire[11:0] T185;
  wire[7:0] T186;
  reg [2:0] acquire_type;
  wire[2:0] T187;
  wire[2:0] T188;
  wire[2:0] T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire[2:0] T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire[25:0] T214;
  wire[25:0] T215;
  wire T216;
  wire T217;
  wire[19:0] T218;
  wire[31:0] T219;
  wire T220;
  wire T221;
  wire T222;
  wire rpq_io_enq_ready;
  wire T223;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_count = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_tag = {1{$random}};
    line_state_state = {1{$random}};
    req_data = {2{$random}};
    acquire_type = {1{$random}};
  end
`endif

  assign T0 = io_mem_finish_ready & can_finish;
  assign can_finish = T63 | T1;
  assign T1 = state == 4'h5;
  assign T2 = reset ? 4'h0 : T3;
  assign T3 = T61 ? T59 : T4;
  assign T4 = T57 ? 4'h4 : T5;
  assign T5 = T35 ? 4'h6 : T6;
  assign T6 = T34 ? 4'h2 : T7;
  assign T7 = T32 ? 4'h3 : T8;
  assign T8 = T30 ? 4'h4 : T9;
  assign T9 = T29 ? 4'h5 : T10;
  assign T10 = T20 ? 4'h6 : T11;
  assign T11 = T18 ? 4'h7 : T12;
  assign T12 = T17 ? 4'h8 : T13;
  assign T13 = T14 ? 4'h0 : state;
  assign T14 = T16 & T15;
  assign T15 = rpq_io_deq_valid ^ 1'h1;
  assign T16 = state == 4'h8;
  assign T17 = state == 4'h7;
  assign T18 = T19 & io_meta_write_ready;
  assign T19 = state == 4'h6;
  assign T20 = T27 & refill_done;
  assign refill_done = reply & T21;
  assign T21 = refill_count == 2'h3;
  assign T22 = T28 ? 2'h0 : T23;
  assign T23 = T25 ? T24 : refill_count;
  assign T24 = refill_count + 2'h1;
  assign T25 = T27 & reply;
  assign reply = io_mem_grant_valid & T26;
  assign T26 = io_mem_grant_bits_payload_client_xact_id == 4'h0;
  assign T27 = state == 4'h5;
  assign T28 = io_req_pri_val & io_req_pri_rdy;
  assign T29 = io_mem_req_ready & io_mem_req_valid;
  assign T30 = T31 & io_meta_write_ready;
  assign T31 = state == 4'h3;
  assign T32 = T33 & reply;
  assign T33 = state == 4'h2;
  assign T34 = io_wb_req_ready & io_wb_req_valid;
  assign T35 = T56 & T36;
  assign T36 = T45 ? T42 : T37;
  assign T37 = T39 | T38;
  assign T38 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T39 = T41 | T40;
  assign T40 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T41 = io_req_bits_old_meta_coh_state == 2'h1;
  assign T42 = T44 | T43;
  assign T43 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T44 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T45 = T47 | T46;
  assign T46 = io_req_bits_cmd == 5'h6;
  assign T47 = T49 | T48;
  assign T48 = io_req_bits_cmd == 5'h3;
  assign T49 = T53 | T50;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h4;
  assign T52 = io_req_bits_cmd[2'h3:2'h3];
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h7;
  assign T55 = io_req_bits_cmd == 5'h1;
  assign T56 = T28 & io_req_bits_tag_match;
  assign T57 = T56 & T58;
  assign T58 = T36 ^ 1'h1;
  assign T59 = T60 ? 4'h1 : 4'h3;
  assign T60 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T61 = T28 & T62;
  assign T62 = io_req_bits_tag_match ^ 1'h1;
  assign T63 = T65 | T64;
  assign T64 = state == 4'h4;
  assign T65 = state == 4'h0;
  assign T66 = T68 & T67;
  assign T67 = io_mem_grant_bits_payload_g_type != 4'h0;
  assign T68 = wb_done | refill_done;
  assign wb_done = reply & T69;
  assign T69 = state == 4'h2;
  assign T70 = T75 ? 1'h0 : T71;
  assign T71 = T73 | T72;
  assign T72 = state == 4'h0;
  assign T73 = io_replay_ready & T74;
  assign T74 = state == 4'h8;
  assign T75 = io_meta_read_ready ^ 1'h1;
  assign T76 = T81 & T77;
  assign T77 = T78 ^ 1'h1;
  assign T78 = T80 | T79;
  assign T79 = io_req_bits_cmd == 5'h3;
  assign T80 = io_req_bits_cmd == 5'h2;
  assign T81 = T128 | T82;
  assign T82 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T83;
  assign T83 = T120 | T84;
  assign T84 = T117 & T85;
  assign T85 = T86 ^ 1'h1;
  assign T86 = T100 | T87;
  assign T87 = T89 & T88;
  assign T88 = io_mem_req_bits_a_type != 3'h1;
  assign T89 = T91 | T90;
  assign T90 = io_req_bits_cmd == 5'h6;
  assign T91 = T93 | T92;
  assign T92 = io_req_bits_cmd == 5'h3;
  assign T93 = T97 | T94;
  assign T94 = T96 | T95;
  assign T95 = io_req_bits_cmd == 5'h4;
  assign T96 = io_req_bits_cmd[2'h3:2'h3];
  assign T97 = T99 | T98;
  assign T98 = io_req_bits_cmd == 5'h7;
  assign T99 = io_req_bits_cmd == 5'h1;
  assign T100 = T110 & T101;
  assign T101 = T103 | T102;
  assign T102 = 3'h6 == io_mem_req_bits_a_type;
  assign T103 = T105 | T104;
  assign T104 = 3'h5 == io_mem_req_bits_a_type;
  assign T105 = T107 | T106;
  assign T106 = 3'h4 == io_mem_req_bits_a_type;
  assign T107 = T109 | T108;
  assign T108 = 3'h3 == io_mem_req_bits_a_type;
  assign T109 = 3'h2 == io_mem_req_bits_a_type;
  assign T110 = T114 | T111;
  assign T111 = T113 | T112;
  assign T112 = io_req_bits_cmd == 5'h4;
  assign T113 = io_req_bits_cmd[2'h3:2'h3];
  assign T114 = T116 | T115;
  assign T115 = io_req_bits_cmd == 5'h6;
  assign T116 = io_req_bits_cmd == 5'h0;
  assign T117 = T119 | T118;
  assign T118 = state == 4'h5;
  assign T119 = state == 4'h4;
  assign T120 = T122 | T121;
  assign T121 = state == 4'h3;
  assign T122 = T124 | T123;
  assign T123 = state == 4'h2;
  assign T124 = state == 4'h1;
  assign idx_match = T126 == T125;
  assign T125 = io_req_bits_addr[4'hb:3'h6];
  assign T126 = req_addr[4'hb:3'h6];
  assign T127 = T28 ? io_req_bits_addr : req_addr;
  assign T128 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T129;
  assign T129 = T143 | T130;
  assign T130 = T138 & T131;
  assign T131 = meta_hazard == 2'h0;
  assign T132 = reset ? 2'h0 : T133;
  assign T133 = T137 ? 2'h1 : T134;
  assign T134 = T136 ? T135 : meta_hazard;
  assign T135 = meta_hazard + 2'h1;
  assign T136 = meta_hazard != 2'h0;
  assign T137 = io_meta_write_ready & io_meta_write_valid;
  assign T138 = T140 & T139;
  assign T139 = state != 4'h3;
  assign T140 = T142 & T141;
  assign T141 = state != 4'h2;
  assign T142 = state != 4'h1;
  assign T143 = idx_match ^ 1'h1;
  assign io_wb_req_bits_r_type = 3'h0;
  assign io_wb_req_bits_master_xact_id = 4'h0;
  assign io_wb_req_bits_client_xact_id = 4'h0;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T144 = T28 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_idx = T126;
  assign io_wb_req_bits_tag = req_old_meta_tag;
  assign T145 = T28 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_valid = T146;
  assign T146 = T147 & ackq_io_enq_ready;
  assign T147 = state == 4'h1;
  assign io_mem_finish_bits_payload_master_xact_id = ackq_io_deq_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = ackq_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ackq_io_deq_bits_header_src;
  assign io_mem_finish_valid = T148;
  assign T148 = ackq_io_deq_valid & can_finish;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_cmd = T149;
  assign T149 = T75 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_data = rpq_io_deq_bits_data;
  assign io_replay_bits_addr = T150;
  assign T150 = {12'h0, T151};
  assign T151 = T152;
  assign T152 = {io_tag, T153};
  assign T153 = {T126, T154};
  assign T154 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_valid = T155;
  assign T155 = T156 & rpq_io_deq_valid;
  assign T156 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T157;
  assign T157 = T158[1'h1:1'h0];
  assign T158 = T178 ? meta_on_flush_state : line_state_state;
  assign T159 = T35 ? meta_on_hit_state : T160;
  assign T160 = T28 ? meta_on_flush_state : T161;
  assign T161 = T25 ? meta_on_grant_state : line_state_state;
  assign meta_on_grant_state = T162;
  assign T162 = T169 ? 2'h1 : T163;
  assign T163 = T168 ? T166 : T164;
  assign T164 = T165 ? 2'h3 : 2'h0;
  assign T165 = io_mem_grant_bits_payload_g_type == 4'h5;
  assign T166 = T167 ? 2'h3 : 2'h2;
  assign T167 = io_mem_req_bits_a_type == 3'h1;
  assign T168 = io_mem_grant_bits_payload_g_type == 4'h2;
  assign T169 = io_mem_grant_bits_payload_g_type == 4'h1;
  assign meta_on_flush_state = 2'h0;
  assign meta_on_hit_state = T170;
  assign T170 = T171 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign T171 = T175 | T172;
  assign T172 = T174 | T173;
  assign T173 = io_req_bits_cmd == 5'h4;
  assign T174 = io_req_bits_cmd[2'h3:2'h3];
  assign T175 = T177 | T176;
  assign T176 = io_req_bits_cmd == 5'h7;
  assign T177 = io_req_bits_cmd == 5'h1;
  assign T178 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = T126;
  assign io_meta_write_valid = T179;
  assign T179 = T181 | T180;
  assign T180 = state == 4'h3;
  assign T181 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = T126;
  assign io_meta_read_valid = T182;
  assign T182 = state == 4'h8;
  assign io_mem_resp_data = T183;
  assign T183 = {64'h0, req_data};
  assign T184 = T28 ? io_req_bits_data : req_data;
  assign io_mem_resp_addr = T185;
  assign T185 = T186 << 3'h4;
  assign T186 = {T126, refill_count};
  assign io_mem_resp_way_en = req_way_en;
  assign io_mem_req_bits_a_type = acquire_type;
  assign T187 = T28 ? T202 : T188;
  assign T188 = T201 ? T189 : acquire_type;
  assign T189 = T190 ? 3'h1 : io_mem_req_bits_a_type;
  assign T190 = T192 | T191;
  assign T191 = io_req_bits_cmd == 5'h6;
  assign T192 = T194 | T193;
  assign T193 = io_req_bits_cmd == 5'h3;
  assign T194 = T198 | T195;
  assign T195 = T197 | T196;
  assign T196 = io_req_bits_cmd == 5'h4;
  assign T197 = io_req_bits_cmd[2'h3:2'h3];
  assign T198 = T200 | T199;
  assign T199 = io_req_bits_cmd == 5'h7;
  assign T200 = io_req_bits_cmd == 5'h1;
  assign T201 = io_req_sec_val & io_req_sec_rdy;
  assign T202 = T203 ? 3'h1 : 3'h0;
  assign T203 = T205 | T204;
  assign T204 = io_req_bits_cmd == 5'h6;
  assign T205 = T207 | T206;
  assign T206 = io_req_bits_cmd == 5'h3;
  assign T207 = T211 | T208;
  assign T208 = T210 | T209;
  assign T209 = io_req_bits_cmd == 5'h4;
  assign T210 = io_req_bits_cmd[2'h3:2'h3];
  assign T211 = T213 | T212;
  assign T212 = io_req_bits_cmd == 5'h7;
  assign T213 = io_req_bits_cmd == 5'h1;
  assign io_mem_req_bits_client_xact_id = 4'h0;
  assign io_mem_req_bits_addr = T214;
  assign T214 = T215;
  assign T215 = {io_tag, T126};
  assign io_mem_req_valid = T216;
  assign T216 = T217 & ackq_io_enq_ready;
  assign T217 = state == 4'h4;
  assign io_tag = T218;
  assign T218 = T219[5'h13:1'h0];
  assign T219 = req_addr >> 4'hc;
  assign io_idx_match = T220;
  assign T220 = T221 & idx_match;
  assign T221 = state != 4'h0;
  assign io_req_sec_rdy = T222;
  assign T222 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T223;
  assign T223 = state == 4'h0;
  Queue_1 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T76 ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_data( io_req_bits_data ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_sdq_id( io_req_sdq_id ),
       .io_deq_ready( T70 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_data( rpq_io_deq_bits_data ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );
  Queue_0 ackq(.clk(clk), .reset(reset),
       .io_enq_ready( ackq_io_enq_ready ),
       .io_enq_valid( T66 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( io_mem_grant_bits_header_src ),
       .io_enq_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_deq_ready( T0 ),
       .io_deq_valid( ackq_io_deq_valid ),
       .io_deq_bits_header_src( ackq_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ackq_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( ackq_io_deq_bits_payload_master_xact_id )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign ackq.io_enq_bits_header_src = {1{$random}};
  `endif

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T61) begin
      state <= T59;
    end else if(T57) begin
      state <= 4'h4;
    end else if(T35) begin
      state <= 4'h6;
    end else if(T34) begin
      state <= 4'h2;
    end else if(T32) begin
      state <= 4'h3;
    end else if(T30) begin
      state <= 4'h4;
    end else if(T29) begin
      state <= 4'h5;
    end else if(T20) begin
      state <= 4'h6;
    end else if(T18) begin
      state <= 4'h7;
    end else if(T17) begin
      state <= 4'h8;
    end else if(T14) begin
      state <= 4'h0;
    end
    if(T28) begin
      refill_count <= 2'h0;
    end else if(T25) begin
      refill_count <= T24;
    end
    if(T28) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T137) begin
      meta_hazard <= 2'h1;
    end else if(T136) begin
      meta_hazard <= T135;
    end
    if(T28) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T28) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(T35) begin
      line_state_state <= meta_on_hit_state;
    end else if(T28) begin
      line_state_state <= meta_on_flush_state;
    end else if(T25) begin
      line_state_state <= meta_on_grant_state;
    end
    if(T28) begin
      req_data <= io_req_bits_data;
    end
    if(T28) begin
      acquire_type <= T202;
    end else if(T201) begin
      acquire_type <= T189;
    end
  end
endmodule

module MSHR_1(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input  io_req_bits_kill,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [63:0] io_req_bits_data,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input  io_req_bits_way_en,
    input [4:0] io_req_sdq_id,
    output io_idx_match,
    output[19:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[3:0] io_mem_req_bits_client_xact_id,
    //output[511:0] io_mem_req_bits_data
    output[2:0] io_mem_req_bits_a_type,
    //output[5:0] io_mem_req_bits_write_mask
    //output[2:0] io_mem_req_bits_subword_addr
    //output[3:0] io_mem_req_bits_atomic_opcode
    output io_mem_resp_way_en,
    output[11:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[127:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[63:0] io_replay_bits_data,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [3:0] io_mem_grant_bits_payload_client_xact_id,
    input [3:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[3:0] io_mem_finish_bits_payload_master_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[19:0] io_wb_req_bits_tag,
    output[5:0] io_wb_req_bits_idx,
    output io_wb_req_bits_way_en,
    output[3:0] io_wb_req_bits_client_xact_id,
    output[3:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy
);

  wire T0;
  wire can_finish;
  wire T1;
  reg [3:0] state;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire rpq_io_deq_valid;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire refill_done;
  wire T21;
  reg [1:0] refill_count;
  wire[1:0] T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire reply;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[3:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire wb_done;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire sec_rdy;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire idx_match;
  wire[5:0] T125;
  wire[5:0] T126;
  reg [43:0] req_addr;
  wire[43:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg [1:0] meta_hazard;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  reg  req_way_en;
  wire T144;
  reg [19:0] req_old_meta_tag;
  wire[19:0] T145;
  wire T146;
  wire ackq_io_enq_ready;
  wire T147;
  wire[3:0] ackq_io_deq_bits_payload_master_xact_id;
  wire[1:0] ackq_io_deq_bits_header_dst;
  wire[1:0] ackq_io_deq_bits_header_src;
  wire T148;
  wire ackq_io_deq_valid;
  wire[4:0] rpq_io_deq_bits_sdq_id;
  wire[4:0] T149;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[7:0] rpq_io_deq_bits_tag;
  wire[63:0] rpq_io_deq_bits_data;
  wire[43:0] T150;
  wire[31:0] T151;
  wire[31:0] T152;
  wire[11:0] T153;
  wire[5:0] T154;
  wire[43:0] rpq_io_deq_bits_addr;
  wire[2:0] rpq_io_deq_bits_typ;
  wire rpq_io_deq_bits_kill;
  wire T155;
  wire T156;
  wire[1:0] T157;
  wire[1:0] T158;
  reg [1:0] line_state_state;
  wire[1:0] T159;
  wire[1:0] T160;
  wire[1:0] T161;
  wire[1:0] meta_on_grant_state;
  wire[1:0] T162;
  wire[1:0] T163;
  wire[1:0] T164;
  wire T165;
  wire[1:0] T166;
  wire T167;
  wire T168;
  wire T169;
  wire[1:0] meta_on_flush_state;
  wire[1:0] meta_on_hit_state;
  wire[1:0] T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire[127:0] T183;
  reg [63:0] req_data;
  wire[63:0] T184;
  wire[11:0] T185;
  wire[7:0] T186;
  reg [2:0] acquire_type;
  wire[2:0] T187;
  wire[2:0] T188;
  wire[2:0] T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire[2:0] T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire[25:0] T214;
  wire[25:0] T215;
  wire T216;
  wire T217;
  wire[19:0] T218;
  wire[31:0] T219;
  wire T220;
  wire T221;
  wire T222;
  wire rpq_io_enq_ready;
  wire T223;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_count = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_tag = {1{$random}};
    line_state_state = {1{$random}};
    req_data = {2{$random}};
    acquire_type = {1{$random}};
  end
`endif

  assign T0 = io_mem_finish_ready & can_finish;
  assign can_finish = T63 | T1;
  assign T1 = state == 4'h5;
  assign T2 = reset ? 4'h0 : T3;
  assign T3 = T61 ? T59 : T4;
  assign T4 = T57 ? 4'h4 : T5;
  assign T5 = T35 ? 4'h6 : T6;
  assign T6 = T34 ? 4'h2 : T7;
  assign T7 = T32 ? 4'h3 : T8;
  assign T8 = T30 ? 4'h4 : T9;
  assign T9 = T29 ? 4'h5 : T10;
  assign T10 = T20 ? 4'h6 : T11;
  assign T11 = T18 ? 4'h7 : T12;
  assign T12 = T17 ? 4'h8 : T13;
  assign T13 = T14 ? 4'h0 : state;
  assign T14 = T16 & T15;
  assign T15 = rpq_io_deq_valid ^ 1'h1;
  assign T16 = state == 4'h8;
  assign T17 = state == 4'h7;
  assign T18 = T19 & io_meta_write_ready;
  assign T19 = state == 4'h6;
  assign T20 = T27 & refill_done;
  assign refill_done = reply & T21;
  assign T21 = refill_count == 2'h3;
  assign T22 = T28 ? 2'h0 : T23;
  assign T23 = T25 ? T24 : refill_count;
  assign T24 = refill_count + 2'h1;
  assign T25 = T27 & reply;
  assign reply = io_mem_grant_valid & T26;
  assign T26 = io_mem_grant_bits_payload_client_xact_id == 4'h1;
  assign T27 = state == 4'h5;
  assign T28 = io_req_pri_val & io_req_pri_rdy;
  assign T29 = io_mem_req_ready & io_mem_req_valid;
  assign T30 = T31 & io_meta_write_ready;
  assign T31 = state == 4'h3;
  assign T32 = T33 & reply;
  assign T33 = state == 4'h2;
  assign T34 = io_wb_req_ready & io_wb_req_valid;
  assign T35 = T56 & T36;
  assign T36 = T45 ? T42 : T37;
  assign T37 = T39 | T38;
  assign T38 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T39 = T41 | T40;
  assign T40 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T41 = io_req_bits_old_meta_coh_state == 2'h1;
  assign T42 = T44 | T43;
  assign T43 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T44 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T45 = T47 | T46;
  assign T46 = io_req_bits_cmd == 5'h6;
  assign T47 = T49 | T48;
  assign T48 = io_req_bits_cmd == 5'h3;
  assign T49 = T53 | T50;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h4;
  assign T52 = io_req_bits_cmd[2'h3:2'h3];
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h7;
  assign T55 = io_req_bits_cmd == 5'h1;
  assign T56 = T28 & io_req_bits_tag_match;
  assign T57 = T56 & T58;
  assign T58 = T36 ^ 1'h1;
  assign T59 = T60 ? 4'h1 : 4'h3;
  assign T60 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T61 = T28 & T62;
  assign T62 = io_req_bits_tag_match ^ 1'h1;
  assign T63 = T65 | T64;
  assign T64 = state == 4'h4;
  assign T65 = state == 4'h0;
  assign T66 = T68 & T67;
  assign T67 = io_mem_grant_bits_payload_g_type != 4'h0;
  assign T68 = wb_done | refill_done;
  assign wb_done = reply & T69;
  assign T69 = state == 4'h2;
  assign T70 = T75 ? 1'h0 : T71;
  assign T71 = T73 | T72;
  assign T72 = state == 4'h0;
  assign T73 = io_replay_ready & T74;
  assign T74 = state == 4'h8;
  assign T75 = io_meta_read_ready ^ 1'h1;
  assign T76 = T81 & T77;
  assign T77 = T78 ^ 1'h1;
  assign T78 = T80 | T79;
  assign T79 = io_req_bits_cmd == 5'h3;
  assign T80 = io_req_bits_cmd == 5'h2;
  assign T81 = T128 | T82;
  assign T82 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T83;
  assign T83 = T120 | T84;
  assign T84 = T117 & T85;
  assign T85 = T86 ^ 1'h1;
  assign T86 = T100 | T87;
  assign T87 = T89 & T88;
  assign T88 = io_mem_req_bits_a_type != 3'h1;
  assign T89 = T91 | T90;
  assign T90 = io_req_bits_cmd == 5'h6;
  assign T91 = T93 | T92;
  assign T92 = io_req_bits_cmd == 5'h3;
  assign T93 = T97 | T94;
  assign T94 = T96 | T95;
  assign T95 = io_req_bits_cmd == 5'h4;
  assign T96 = io_req_bits_cmd[2'h3:2'h3];
  assign T97 = T99 | T98;
  assign T98 = io_req_bits_cmd == 5'h7;
  assign T99 = io_req_bits_cmd == 5'h1;
  assign T100 = T110 & T101;
  assign T101 = T103 | T102;
  assign T102 = 3'h6 == io_mem_req_bits_a_type;
  assign T103 = T105 | T104;
  assign T104 = 3'h5 == io_mem_req_bits_a_type;
  assign T105 = T107 | T106;
  assign T106 = 3'h4 == io_mem_req_bits_a_type;
  assign T107 = T109 | T108;
  assign T108 = 3'h3 == io_mem_req_bits_a_type;
  assign T109 = 3'h2 == io_mem_req_bits_a_type;
  assign T110 = T114 | T111;
  assign T111 = T113 | T112;
  assign T112 = io_req_bits_cmd == 5'h4;
  assign T113 = io_req_bits_cmd[2'h3:2'h3];
  assign T114 = T116 | T115;
  assign T115 = io_req_bits_cmd == 5'h6;
  assign T116 = io_req_bits_cmd == 5'h0;
  assign T117 = T119 | T118;
  assign T118 = state == 4'h5;
  assign T119 = state == 4'h4;
  assign T120 = T122 | T121;
  assign T121 = state == 4'h3;
  assign T122 = T124 | T123;
  assign T123 = state == 4'h2;
  assign T124 = state == 4'h1;
  assign idx_match = T126 == T125;
  assign T125 = io_req_bits_addr[4'hb:3'h6];
  assign T126 = req_addr[4'hb:3'h6];
  assign T127 = T28 ? io_req_bits_addr : req_addr;
  assign T128 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T129;
  assign T129 = T143 | T130;
  assign T130 = T138 & T131;
  assign T131 = meta_hazard == 2'h0;
  assign T132 = reset ? 2'h0 : T133;
  assign T133 = T137 ? 2'h1 : T134;
  assign T134 = T136 ? T135 : meta_hazard;
  assign T135 = meta_hazard + 2'h1;
  assign T136 = meta_hazard != 2'h0;
  assign T137 = io_meta_write_ready & io_meta_write_valid;
  assign T138 = T140 & T139;
  assign T139 = state != 4'h3;
  assign T140 = T142 & T141;
  assign T141 = state != 4'h2;
  assign T142 = state != 4'h1;
  assign T143 = idx_match ^ 1'h1;
  assign io_wb_req_bits_r_type = 3'h0;
  assign io_wb_req_bits_master_xact_id = 4'h0;
  assign io_wb_req_bits_client_xact_id = 4'h1;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T144 = T28 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_idx = T126;
  assign io_wb_req_bits_tag = req_old_meta_tag;
  assign T145 = T28 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_valid = T146;
  assign T146 = T147 & ackq_io_enq_ready;
  assign T147 = state == 4'h1;
  assign io_mem_finish_bits_payload_master_xact_id = ackq_io_deq_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = ackq_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ackq_io_deq_bits_header_src;
  assign io_mem_finish_valid = T148;
  assign T148 = ackq_io_deq_valid & can_finish;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_cmd = T149;
  assign T149 = T75 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_data = rpq_io_deq_bits_data;
  assign io_replay_bits_addr = T150;
  assign T150 = {12'h0, T151};
  assign T151 = T152;
  assign T152 = {io_tag, T153};
  assign T153 = {T126, T154};
  assign T154 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_valid = T155;
  assign T155 = T156 & rpq_io_deq_valid;
  assign T156 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T157;
  assign T157 = T158[1'h1:1'h0];
  assign T158 = T178 ? meta_on_flush_state : line_state_state;
  assign T159 = T35 ? meta_on_hit_state : T160;
  assign T160 = T28 ? meta_on_flush_state : T161;
  assign T161 = T25 ? meta_on_grant_state : line_state_state;
  assign meta_on_grant_state = T162;
  assign T162 = T169 ? 2'h1 : T163;
  assign T163 = T168 ? T166 : T164;
  assign T164 = T165 ? 2'h3 : 2'h0;
  assign T165 = io_mem_grant_bits_payload_g_type == 4'h5;
  assign T166 = T167 ? 2'h3 : 2'h2;
  assign T167 = io_mem_req_bits_a_type == 3'h1;
  assign T168 = io_mem_grant_bits_payload_g_type == 4'h2;
  assign T169 = io_mem_grant_bits_payload_g_type == 4'h1;
  assign meta_on_flush_state = 2'h0;
  assign meta_on_hit_state = T170;
  assign T170 = T171 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign T171 = T175 | T172;
  assign T172 = T174 | T173;
  assign T173 = io_req_bits_cmd == 5'h4;
  assign T174 = io_req_bits_cmd[2'h3:2'h3];
  assign T175 = T177 | T176;
  assign T176 = io_req_bits_cmd == 5'h7;
  assign T177 = io_req_bits_cmd == 5'h1;
  assign T178 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = T126;
  assign io_meta_write_valid = T179;
  assign T179 = T181 | T180;
  assign T180 = state == 4'h3;
  assign T181 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = T126;
  assign io_meta_read_valid = T182;
  assign T182 = state == 4'h8;
  assign io_mem_resp_data = T183;
  assign T183 = {64'h0, req_data};
  assign T184 = T28 ? io_req_bits_data : req_data;
  assign io_mem_resp_addr = T185;
  assign T185 = T186 << 3'h4;
  assign T186 = {T126, refill_count};
  assign io_mem_resp_way_en = req_way_en;
  assign io_mem_req_bits_a_type = acquire_type;
  assign T187 = T28 ? T202 : T188;
  assign T188 = T201 ? T189 : acquire_type;
  assign T189 = T190 ? 3'h1 : io_mem_req_bits_a_type;
  assign T190 = T192 | T191;
  assign T191 = io_req_bits_cmd == 5'h6;
  assign T192 = T194 | T193;
  assign T193 = io_req_bits_cmd == 5'h3;
  assign T194 = T198 | T195;
  assign T195 = T197 | T196;
  assign T196 = io_req_bits_cmd == 5'h4;
  assign T197 = io_req_bits_cmd[2'h3:2'h3];
  assign T198 = T200 | T199;
  assign T199 = io_req_bits_cmd == 5'h7;
  assign T200 = io_req_bits_cmd == 5'h1;
  assign T201 = io_req_sec_val & io_req_sec_rdy;
  assign T202 = T203 ? 3'h1 : 3'h0;
  assign T203 = T205 | T204;
  assign T204 = io_req_bits_cmd == 5'h6;
  assign T205 = T207 | T206;
  assign T206 = io_req_bits_cmd == 5'h3;
  assign T207 = T211 | T208;
  assign T208 = T210 | T209;
  assign T209 = io_req_bits_cmd == 5'h4;
  assign T210 = io_req_bits_cmd[2'h3:2'h3];
  assign T211 = T213 | T212;
  assign T212 = io_req_bits_cmd == 5'h7;
  assign T213 = io_req_bits_cmd == 5'h1;
  assign io_mem_req_bits_client_xact_id = 4'h1;
  assign io_mem_req_bits_addr = T214;
  assign T214 = T215;
  assign T215 = {io_tag, T126};
  assign io_mem_req_valid = T216;
  assign T216 = T217 & ackq_io_enq_ready;
  assign T217 = state == 4'h4;
  assign io_tag = T218;
  assign T218 = T219[5'h13:1'h0];
  assign T219 = req_addr >> 4'hc;
  assign io_idx_match = T220;
  assign T220 = T221 & idx_match;
  assign T221 = state != 4'h0;
  assign io_req_sec_rdy = T222;
  assign T222 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T223;
  assign T223 = state == 4'h0;
  Queue_1 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T76 ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_data( io_req_bits_data ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_sdq_id( io_req_sdq_id ),
       .io_deq_ready( T70 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_data( rpq_io_deq_bits_data ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );
  Queue_0 ackq(.clk(clk), .reset(reset),
       .io_enq_ready( ackq_io_enq_ready ),
       .io_enq_valid( T66 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( io_mem_grant_bits_header_src ),
       .io_enq_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_deq_ready( T0 ),
       .io_deq_valid( ackq_io_deq_valid ),
       .io_deq_bits_header_src( ackq_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ackq_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( ackq_io_deq_bits_payload_master_xact_id )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign ackq.io_enq_bits_header_src = {1{$random}};
  `endif

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T61) begin
      state <= T59;
    end else if(T57) begin
      state <= 4'h4;
    end else if(T35) begin
      state <= 4'h6;
    end else if(T34) begin
      state <= 4'h2;
    end else if(T32) begin
      state <= 4'h3;
    end else if(T30) begin
      state <= 4'h4;
    end else if(T29) begin
      state <= 4'h5;
    end else if(T20) begin
      state <= 4'h6;
    end else if(T18) begin
      state <= 4'h7;
    end else if(T17) begin
      state <= 4'h8;
    end else if(T14) begin
      state <= 4'h0;
    end
    if(T28) begin
      refill_count <= 2'h0;
    end else if(T25) begin
      refill_count <= T24;
    end
    if(T28) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T137) begin
      meta_hazard <= 2'h1;
    end else if(T136) begin
      meta_hazard <= T135;
    end
    if(T28) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T28) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(T35) begin
      line_state_state <= meta_on_hit_state;
    end else if(T28) begin
      line_state_state <= meta_on_flush_state;
    end else if(T25) begin
      line_state_state <= meta_on_grant_state;
    end
    if(T28) begin
      req_data <= io_req_bits_data;
    end
    if(T28) begin
      acquire_type <= T202;
    end else if(T201) begin
      acquire_type <= T189;
    end
  end
endmodule

module MSHRFile(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input  io_req_bits_kill,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [63:0] io_req_bits_data,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input  io_req_bits_way_en,
    output io_secondary_miss,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[3:0] io_mem_req_bits_client_xact_id,
    output[511:0] io_mem_req_bits_data,
    output[2:0] io_mem_req_bits_a_type,
    output[5:0] io_mem_req_bits_write_mask,
    output[2:0] io_mem_req_bits_subword_addr,
    output[3:0] io_mem_req_bits_atomic_opcode,
    output io_mem_resp_way_en,
    output[11:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[127:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[63:0] io_replay_bits_data,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [3:0] io_mem_grant_bits_payload_client_xact_id,
    input [3:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[3:0] io_mem_finish_bits_payload_master_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[19:0] io_wb_req_bits_tag,
    output[5:0] io_wb_req_bits_idx,
    output io_wb_req_bits_way_en,
    output[3:0] io_wb_req_bits_client_xact_id,
    output[3:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy,
    output io_fence_rdy
);

  wire wb_req_arb_io_in_1_ready;
  wire mem_finish_arb_io_in_1_ready;
  wire replay_arb_io_in_1_ready;
  wire meta_write_arb_io_in_1_ready;
  wire meta_read_arb_io_in_1_ready;
  wire mem_req_arb_io_in_1_ready;
  wire[4:0] T0;
  wire[4:0] T1;
  wire[4:0] T2;
  wire[4:0] T3;
  wire[4:0] T4;
  wire[4:0] T5;
  wire[4:0] T6;
  wire[4:0] T7;
  wire[4:0] T8;
  wire[4:0] T9;
  wire[4:0] T10;
  wire[4:0] T11;
  wire[4:0] T12;
  wire[4:0] T13;
  wire[4:0] T14;
  wire[4:0] T15;
  wire T16;
  wire[16:0] T17;
  wire[16:0] T18;
  reg [16:0] sdq_val;
  wire[16:0] T19;
  wire[31:0] T20;
  wire[31:0] T21;
  wire[31:0] T22;
  wire[31:0] T23;
  wire[31:0] T24;
  wire[16:0] T25;
  wire[16:0] T26;
  wire[16:0] T27;
  wire sdq_enq;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[16:0] T36;
  wire[16:0] T37;
  wire[16:0] T38;
  wire[16:0] T39;
  wire[16:0] T40;
  wire[16:0] T41;
  wire[16:0] T42;
  wire[16:0] T43;
  wire[16:0] T44;
  wire[16:0] T45;
  wire[16:0] T46;
  wire[16:0] T47;
  wire[16:0] T48;
  wire[16:0] T49;
  wire[16:0] T50;
  wire[16:0] T51;
  wire[16:0] T52;
  wire T53;
  wire[16:0] T54;
  wire[16:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[31:0] T72;
  wire[31:0] T73;
  wire[31:0] T74;
  wire[31:0] T75;
  wire[16:0] T76;
  wire[16:0] T77;
  wire free_sdq;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire[31:0] T86;
  wire[31:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire tag_match;
  wire[31:0] T105;
  wire[31:0] T106;
  wire[19:0] T107;
  wire[19:0] T108;
  wire[19:0] tagList_1;
  wire[19:0] MSHR_1_io_tag;
  wire idxMatch_1;
  wire MSHR_1_io_idx_match;
  wire[19:0] T109;
  wire[19:0] tagList_0;
  wire[19:0] MSHR_0_io_tag;
  wire idxMatch_0;
  wire MSHR_0_io_idx_match;
  wire T110;
  wire sdq_rdy;
  wire T111;
  wire alloc_arb_io_in_1_ready;
  wire wb_req_arb_io_in_0_ready;
  wire mem_finish_arb_io_in_0_ready;
  wire replay_arb_io_in_0_ready;
  wire meta_write_arb_io_in_0_ready;
  wire meta_read_arb_io_in_0_ready;
  wire mem_req_arb_io_in_0_ready;
  wire T112;
  wire T113;
  wire alloc_arb_io_in_0_ready;
  wire T114;
  wire T115;
  wire idx_match;
  wire T116;
  wire MSHR_0_io_req_pri_rdy;
  wire MSHR_1_io_req_pri_rdy;
  wire[4:0] MSHR_0_io_replay_bits_sdq_id;
  wire[4:0] MSHR_0_io_replay_bits_cmd;
  wire[7:0] MSHR_0_io_replay_bits_tag;
  wire[63:0] MSHR_0_io_replay_bits_data;
  wire[43:0] MSHR_0_io_replay_bits_addr;
  wire MSHR_0_io_replay_bits_phys;
  wire[2:0] MSHR_0_io_replay_bits_typ;
  wire MSHR_0_io_replay_bits_kill;
  wire MSHR_0_io_replay_valid;
  wire[4:0] MSHR_1_io_replay_bits_sdq_id;
  wire[4:0] MSHR_1_io_replay_bits_cmd;
  wire[7:0] MSHR_1_io_replay_bits_tag;
  wire[63:0] MSHR_1_io_replay_bits_data;
  wire[43:0] MSHR_1_io_replay_bits_addr;
  wire MSHR_1_io_replay_bits_phys;
  wire[2:0] MSHR_1_io_replay_bits_typ;
  wire MSHR_1_io_replay_bits_kill;
  wire MSHR_1_io_replay_valid;
  wire[2:0] MSHR_0_io_wb_req_bits_r_type;
  wire[3:0] MSHR_0_io_wb_req_bits_master_xact_id;
  wire[3:0] MSHR_0_io_wb_req_bits_client_xact_id;
  wire MSHR_0_io_wb_req_bits_way_en;
  wire[5:0] MSHR_0_io_wb_req_bits_idx;
  wire[19:0] MSHR_0_io_wb_req_bits_tag;
  wire MSHR_0_io_wb_req_valid;
  wire[2:0] MSHR_1_io_wb_req_bits_r_type;
  wire[3:0] MSHR_1_io_wb_req_bits_master_xact_id;
  wire[3:0] MSHR_1_io_wb_req_bits_client_xact_id;
  wire MSHR_1_io_wb_req_bits_way_en;
  wire[5:0] MSHR_1_io_wb_req_bits_idx;
  wire[19:0] MSHR_1_io_wb_req_bits_tag;
  wire MSHR_1_io_wb_req_valid;
  wire[3:0] MSHR_0_io_mem_finish_bits_payload_master_xact_id;
  wire[1:0] MSHR_0_io_mem_finish_bits_header_dst;
  wire[1:0] MSHR_0_io_mem_finish_bits_header_src;
  wire MSHR_0_io_mem_finish_valid;
  wire[3:0] MSHR_1_io_mem_finish_bits_payload_master_xact_id;
  wire[1:0] MSHR_1_io_mem_finish_bits_header_dst;
  wire[1:0] MSHR_1_io_mem_finish_bits_header_src;
  wire MSHR_1_io_mem_finish_valid;
  wire[2:0] MSHR_0_io_mem_req_bits_a_type;
  wire[3:0] MSHR_0_io_mem_req_bits_client_xact_id;
  wire[25:0] MSHR_0_io_mem_req_bits_addr;
  wire MSHR_0_io_mem_req_valid;
  wire[2:0] MSHR_1_io_mem_req_bits_a_type;
  wire[3:0] MSHR_1_io_mem_req_bits_client_xact_id;
  wire[25:0] MSHR_1_io_mem_req_bits_addr;
  wire MSHR_1_io_mem_req_valid;
  wire[1:0] MSHR_0_io_meta_write_bits_data_coh_state;
  wire[19:0] MSHR_0_io_meta_write_bits_data_tag;
  wire MSHR_0_io_meta_write_bits_way_en;
  wire[5:0] MSHR_0_io_meta_write_bits_idx;
  wire MSHR_0_io_meta_write_valid;
  wire[1:0] MSHR_1_io_meta_write_bits_data_coh_state;
  wire[19:0] MSHR_1_io_meta_write_bits_data_tag;
  wire MSHR_1_io_meta_write_bits_way_en;
  wire[5:0] MSHR_1_io_meta_write_bits_idx;
  wire MSHR_1_io_meta_write_valid;
  wire[19:0] MSHR_0_io_meta_read_bits_tag;
  wire[5:0] MSHR_0_io_meta_read_bits_idx;
  wire MSHR_0_io_meta_read_valid;
  wire[19:0] MSHR_1_io_meta_read_bits_tag;
  wire[5:0] MSHR_1_io_meta_read_bits_idx;
  wire MSHR_1_io_meta_read_valid;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire MSHR_0_io_probe_rdy;
  wire T124;
  wire MSHR_1_io_probe_rdy;
  wire[2:0] wb_req_arb_io_out_bits_r_type;
  wire[3:0] wb_req_arb_io_out_bits_master_xact_id;
  wire[3:0] wb_req_arb_io_out_bits_client_xact_id;
  wire wb_req_arb_io_out_bits_way_en;
  wire[5:0] wb_req_arb_io_out_bits_idx;
  wire[19:0] wb_req_arb_io_out_bits_tag;
  wire wb_req_arb_io_out_valid;
  wire[3:0] mem_finish_arb_io_out_bits_payload_master_xact_id;
  wire[1:0] mem_finish_arb_io_out_bits_header_dst;
  wire[1:0] mem_finish_arb_io_out_bits_header_src;
  wire mem_finish_arb_io_out_valid;
  wire[4:0] replay_arb_io_out_bits_sdq_id;
  wire[4:0] replay_arb_io_out_bits_cmd;
  wire[7:0] replay_arb_io_out_bits_tag;
  wire[63:0] T125;
  reg [63:0] sdq [16:0];
  wire[63:0] T126;
  wire T127;
  wire T128;
  wire[4:0] T129;
  reg [4:0] R130;
  wire[4:0] T131;
  wire[43:0] replay_arb_io_out_bits_addr;
  wire replay_arb_io_out_bits_phys;
  wire[2:0] replay_arb_io_out_bits_typ;
  wire replay_arb_io_out_bits_kill;
  wire replay_arb_io_out_valid;
  wire[1:0] meta_write_arb_io_out_bits_data_coh_state;
  wire[19:0] meta_write_arb_io_out_bits_data_tag;
  wire meta_write_arb_io_out_bits_way_en;
  wire[5:0] meta_write_arb_io_out_bits_idx;
  wire meta_write_arb_io_out_valid;
  wire[19:0] meta_read_arb_io_out_bits_tag;
  wire[5:0] meta_read_arb_io_out_bits_idx;
  wire meta_read_arb_io_out_valid;
  wire[127:0] T132;
  wire[127:0] memRespMux_0_data;
  wire[127:0] MSHR_0_io_mem_resp_data;
  wire[127:0] memRespMux_1_data;
  wire[127:0] MSHR_1_io_mem_resp_data;
  wire T133;
  wire T134;
  wire[1:0] T135;
  wire[1:0] memRespMux_0_wmask;
  wire[1:0] MSHR_0_io_mem_resp_wmask;
  wire[1:0] memRespMux_1_wmask;
  wire[1:0] MSHR_1_io_mem_resp_wmask;
  wire[11:0] T136;
  wire[11:0] memRespMux_0_addr;
  wire[11:0] MSHR_0_io_mem_resp_addr;
  wire[11:0] memRespMux_1_addr;
  wire[11:0] MSHR_1_io_mem_resp_addr;
  wire T137;
  wire memRespMux_0_way_en;
  wire MSHR_0_io_mem_resp_way_en;
  wire memRespMux_1_way_en;
  wire MSHR_1_io_mem_resp_way_en;
  wire[3:0] mem_req_arb_io_out_bits_atomic_opcode;
  wire[2:0] mem_req_arb_io_out_bits_subword_addr;
  wire[5:0] mem_req_arb_io_out_bits_write_mask;
  wire[2:0] mem_req_arb_io_out_bits_a_type;
  wire[511:0] mem_req_arb_io_out_bits_data;
  wire[3:0] mem_req_arb_io_out_bits_client_xact_id;
  wire[25:0] mem_req_arb_io_out_bits_addr;
  wire mem_req_arb_io_out_valid;
  wire T138;
  wire T139;
  wire pri_rdy;
  wire T140;
  wire sec_rdy;
  wire MSHR_1_io_req_sec_rdy;
  wire MSHR_0_io_req_sec_rdy;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    sdq_val = {1{$random}};
    for (initvar = 0; initvar < 17; initvar = initvar+1)
      sdq[initvar] = {2{$random}};
    R130 = {1{$random}};
  end
`endif

  assign T0 = T103 ? 1'h0 : T1;
  assign T1 = T102 ? 1'h1 : T2;
  assign T2 = T101 ? 2'h2 : T3;
  assign T3 = T100 ? 2'h3 : T4;
  assign T4 = T99 ? 3'h4 : T5;
  assign T5 = T98 ? 3'h5 : T6;
  assign T6 = T97 ? 3'h6 : T7;
  assign T7 = T96 ? 3'h7 : T8;
  assign T8 = T95 ? 4'h8 : T9;
  assign T9 = T94 ? 4'h9 : T10;
  assign T10 = T93 ? 4'ha : T11;
  assign T11 = T92 ? 4'hb : T12;
  assign T12 = T91 ? 4'hc : T13;
  assign T13 = T90 ? 4'hd : T14;
  assign T14 = T89 ? 4'he : T15;
  assign T15 = T16 ? 4'hf : 5'h10;
  assign T16 = T17[4'hf:4'hf];
  assign T17 = ~ T18;
  assign T18 = sdq_val[5'h10:1'h0];
  assign T19 = T20[5'h10:1'h0];
  assign T20 = reset ? 32'h0 : T21;
  assign T21 = T88 ? T23 : T22;
  assign T22 = {15'h0, sdq_val};
  assign T23 = T72 | T24;
  assign T24 = {15'h0, T25};
  assign T25 = T36 & T26;
  assign T26 = 17'h0 - T27;
  assign T27 = {16'h0, sdq_enq};
  assign sdq_enq = T35 & T28;
  assign T28 = T32 | T29;
  assign T29 = T31 | T30;
  assign T30 = io_req_bits_cmd == 5'h4;
  assign T31 = io_req_bits_cmd[2'h3:2'h3];
  assign T32 = T34 | T33;
  assign T33 = io_req_bits_cmd == 5'h7;
  assign T34 = io_req_bits_cmd == 5'h1;
  assign T35 = io_req_valid & io_req_ready;
  assign T36 = T71 ? 17'h1 : T37;
  assign T37 = T70 ? 17'h2 : T38;
  assign T38 = T69 ? 17'h4 : T39;
  assign T39 = T68 ? 17'h8 : T40;
  assign T40 = T67 ? 17'h10 : T41;
  assign T41 = T66 ? 17'h20 : T42;
  assign T42 = T65 ? 17'h40 : T43;
  assign T43 = T64 ? 17'h80 : T44;
  assign T44 = T63 ? 17'h100 : T45;
  assign T45 = T62 ? 17'h200 : T46;
  assign T46 = T61 ? 17'h400 : T47;
  assign T47 = T60 ? 17'h800 : T48;
  assign T48 = T59 ? 17'h1000 : T49;
  assign T49 = T58 ? 17'h2000 : T50;
  assign T50 = T57 ? 17'h4000 : T51;
  assign T51 = T56 ? 17'h8000 : T52;
  assign T52 = T53 ? 17'h10000 : 17'h0;
  assign T53 = T54[5'h10:5'h10];
  assign T54 = ~ T55;
  assign T55 = sdq_val[5'h10:1'h0];
  assign T56 = T54[4'hf:4'hf];
  assign T57 = T54[4'he:4'he];
  assign T58 = T54[4'hd:4'hd];
  assign T59 = T54[4'hc:4'hc];
  assign T60 = T54[4'hb:4'hb];
  assign T61 = T54[4'ha:4'ha];
  assign T62 = T54[4'h9:4'h9];
  assign T63 = T54[4'h8:4'h8];
  assign T64 = T54[3'h7:3'h7];
  assign T65 = T54[3'h6:3'h6];
  assign T66 = T54[3'h5:3'h5];
  assign T67 = T54[3'h4:3'h4];
  assign T68 = T54[2'h3:2'h3];
  assign T69 = T54[2'h2:2'h2];
  assign T70 = T54[1'h1:1'h1];
  assign T71 = T54[1'h0:1'h0];
  assign T72 = T87 & T73;
  assign T73 = ~ T74;
  assign T74 = T86 & T75;
  assign T75 = {15'h0, T76};
  assign T76 = 17'h0 - T77;
  assign T77 = {16'h0, free_sdq};
  assign free_sdq = T85 & T78;
  assign T78 = T82 | T79;
  assign T79 = T81 | T80;
  assign T80 = io_replay_bits_cmd == 5'h4;
  assign T81 = io_replay_bits_cmd[2'h3:2'h3];
  assign T82 = T84 | T83;
  assign T83 = io_replay_bits_cmd == 5'h7;
  assign T84 = io_replay_bits_cmd == 5'h1;
  assign T85 = io_replay_ready & io_replay_valid;
  assign T86 = 1'h1 << io_replay_bits_sdq_id;
  assign T87 = {15'h0, sdq_val};
  assign T88 = io_replay_valid | sdq_enq;
  assign T89 = T17[4'he:4'he];
  assign T90 = T17[4'hd:4'hd];
  assign T91 = T17[4'hc:4'hc];
  assign T92 = T17[4'hb:4'hb];
  assign T93 = T17[4'ha:4'ha];
  assign T94 = T17[4'h9:4'h9];
  assign T95 = T17[4'h8:4'h8];
  assign T96 = T17[3'h7:3'h7];
  assign T97 = T17[3'h6:3'h6];
  assign T98 = T17[3'h5:3'h5];
  assign T99 = T17[3'h4:3'h4];
  assign T100 = T17[2'h3:2'h3];
  assign T101 = T17[2'h2:2'h2];
  assign T102 = T17[1'h1:1'h1];
  assign T103 = T17[1'h0:1'h0];
  assign T104 = T110 & tag_match;
  assign tag_match = T106 == T105;
  assign T105 = io_req_bits_addr >> 4'hc;
  assign T106 = {12'h0, T107};
  assign T107 = T109 | T108;
  assign T108 = idxMatch_1 ? tagList_1 : 20'h0;
  assign tagList_1 = MSHR_1_io_tag;
  assign idxMatch_1 = MSHR_1_io_idx_match;
  assign T109 = idxMatch_0 ? tagList_0 : 20'h0;
  assign tagList_0 = MSHR_0_io_tag;
  assign idxMatch_0 = MSHR_0_io_idx_match;
  assign T110 = io_req_valid & sdq_rdy;
  assign sdq_rdy = T111 ^ 1'h1;
  assign T111 = sdq_val == 17'h1ffff;
  assign T112 = T113 & tag_match;
  assign T113 = io_req_valid & sdq_rdy;
  assign T114 = T116 & T115;
  assign T115 = idx_match ^ 1'h1;
  assign idx_match = MSHR_0_io_idx_match | MSHR_1_io_idx_match;
  assign T116 = io_req_valid & sdq_rdy;
  assign io_fence_rdy = T117;
  assign T117 = T120 ? 1'h0 : T118;
  assign T118 = T119 == 1'h0;
  assign T119 = MSHR_0_io_req_pri_rdy ^ 1'h1;
  assign T120 = MSHR_1_io_req_pri_rdy ^ 1'h1;
  assign io_probe_rdy = T121;
  assign T121 = T124 ? 1'h0 : T122;
  assign T122 = T123 == 1'h0;
  assign T123 = MSHR_0_io_probe_rdy ^ 1'h1;
  assign T124 = MSHR_1_io_probe_rdy ^ 1'h1;
  assign io_wb_req_bits_r_type = wb_req_arb_io_out_bits_r_type;
  assign io_wb_req_bits_master_xact_id = wb_req_arb_io_out_bits_master_xact_id;
  assign io_wb_req_bits_client_xact_id = wb_req_arb_io_out_bits_client_xact_id;
  assign io_wb_req_bits_way_en = wb_req_arb_io_out_bits_way_en;
  assign io_wb_req_bits_idx = wb_req_arb_io_out_bits_idx;
  assign io_wb_req_bits_tag = wb_req_arb_io_out_bits_tag;
  assign io_wb_req_valid = wb_req_arb_io_out_valid;
  assign io_mem_finish_bits_payload_master_xact_id = mem_finish_arb_io_out_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = mem_finish_arb_io_out_bits_header_dst;
  assign io_mem_finish_bits_header_src = mem_finish_arb_io_out_bits_header_src;
  assign io_mem_finish_valid = mem_finish_arb_io_out_valid;
  assign io_replay_bits_sdq_id = replay_arb_io_out_bits_sdq_id;
  assign io_replay_bits_cmd = replay_arb_io_out_bits_cmd;
  assign io_replay_bits_tag = replay_arb_io_out_bits_tag;
  assign io_replay_bits_data = T125;
  assign T125 = sdq[R130];
  always @(posedge clk)
    if (T127)
      sdq[T0] <= io_req_bits_data;
  assign T127 = sdq_enq & T128;
  assign T128 = T129 < 5'h11;
  assign T129 = T0[3'h4:1'h0];
  assign T131 = free_sdq ? replay_arb_io_out_bits_sdq_id : R130;
  assign io_replay_bits_addr = replay_arb_io_out_bits_addr;
  assign io_replay_bits_phys = replay_arb_io_out_bits_phys;
  assign io_replay_bits_typ = replay_arb_io_out_bits_typ;
  assign io_replay_bits_kill = replay_arb_io_out_bits_kill;
  assign io_replay_valid = replay_arb_io_out_valid;
  assign io_meta_write_bits_data_coh_state = meta_write_arb_io_out_bits_data_coh_state;
  assign io_meta_write_bits_data_tag = meta_write_arb_io_out_bits_data_tag;
  assign io_meta_write_bits_way_en = meta_write_arb_io_out_bits_way_en;
  assign io_meta_write_bits_idx = meta_write_arb_io_out_bits_idx;
  assign io_meta_write_valid = meta_write_arb_io_out_valid;
  assign io_meta_read_bits_tag = meta_read_arb_io_out_bits_tag;
  assign io_meta_read_bits_idx = meta_read_arb_io_out_bits_idx;
  assign io_meta_read_valid = meta_read_arb_io_out_valid;
  assign io_mem_resp_data = T132;
  assign T132 = T133 ? memRespMux_1_data : memRespMux_0_data;
  assign memRespMux_0_data = MSHR_0_io_mem_resp_data;
  assign memRespMux_1_data = MSHR_1_io_mem_resp_data;
  assign T133 = T134;
  assign T134 = io_mem_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign io_mem_resp_wmask = T135;
  assign T135 = T133 ? memRespMux_1_wmask : memRespMux_0_wmask;
  assign memRespMux_0_wmask = MSHR_0_io_mem_resp_wmask;
  assign memRespMux_1_wmask = MSHR_1_io_mem_resp_wmask;
  assign io_mem_resp_addr = T136;
  assign T136 = T133 ? memRespMux_1_addr : memRespMux_0_addr;
  assign memRespMux_0_addr = MSHR_0_io_mem_resp_addr;
  assign memRespMux_1_addr = MSHR_1_io_mem_resp_addr;
  assign io_mem_resp_way_en = T137;
  assign T137 = T133 ? memRespMux_1_way_en : memRespMux_0_way_en;
  assign memRespMux_0_way_en = MSHR_0_io_mem_resp_way_en;
  assign memRespMux_1_way_en = MSHR_1_io_mem_resp_way_en;
  assign io_mem_req_bits_atomic_opcode = mem_req_arb_io_out_bits_atomic_opcode;
  assign io_mem_req_bits_subword_addr = mem_req_arb_io_out_bits_subword_addr;
  assign io_mem_req_bits_write_mask = mem_req_arb_io_out_bits_write_mask;
  assign io_mem_req_bits_a_type = mem_req_arb_io_out_bits_a_type;
  assign io_mem_req_bits_data = mem_req_arb_io_out_bits_data;
  assign io_mem_req_bits_client_xact_id = mem_req_arb_io_out_bits_client_xact_id;
  assign io_mem_req_bits_addr = mem_req_arb_io_out_bits_addr;
  assign io_mem_req_valid = mem_req_arb_io_out_valid;
  assign io_secondary_miss = idx_match;
  assign io_req_ready = T138;
  assign T138 = T139 & sdq_rdy;
  assign T139 = idx_match ? T140 : pri_rdy;
  assign pri_rdy = MSHR_0_io_req_pri_rdy | MSHR_1_io_req_pri_rdy;
  assign T140 = tag_match & sec_rdy;
  assign sec_rdy = MSHR_0_io_req_sec_rdy | MSHR_1_io_req_sec_rdy;
  Arbiter_0 meta_read_arb(
       .io_in_1_ready( meta_read_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_read_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_in_1_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_in_0_ready( meta_read_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_meta_read_valid ),
       .io_in_0_bits_idx( MSHR_0_io_meta_read_bits_idx ),
       .io_in_0_bits_tag( MSHR_0_io_meta_read_bits_tag ),
       .io_out_ready( io_meta_read_ready ),
       .io_out_valid( meta_read_arb_io_out_valid ),
       .io_out_bits_idx( meta_read_arb_io_out_bits_idx ),
       .io_out_bits_tag( meta_read_arb_io_out_bits_tag )
       //.io_chosen(  )
  );
  Arbiter_1 meta_write_arb(
       .io_in_1_ready( meta_write_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_write_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( meta_write_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_meta_write_valid ),
       .io_in_0_bits_idx( MSHR_0_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( MSHR_0_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( MSHR_0_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( MSHR_0_io_meta_write_bits_data_coh_state ),
       .io_out_ready( io_meta_write_ready ),
       .io_out_valid( meta_write_arb_io_out_valid ),
       .io_out_bits_idx( meta_write_arb_io_out_bits_idx ),
       .io_out_bits_way_en( meta_write_arb_io_out_bits_way_en ),
       .io_out_bits_data_tag( meta_write_arb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( meta_write_arb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  Arbiter_2 mem_req_arb(
       .io_in_1_ready( mem_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_req_valid ),
       .io_in_1_bits_addr( MSHR_1_io_mem_req_bits_addr ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       //.io_in_1_bits_data(  )
       .io_in_1_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       //.io_in_1_bits_write_mask(  )
       //.io_in_1_bits_subword_addr(  )
       //.io_in_1_bits_atomic_opcode(  )
       .io_in_0_ready( mem_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_mem_req_valid ),
       .io_in_0_bits_addr( MSHR_0_io_mem_req_bits_addr ),
       .io_in_0_bits_client_xact_id( MSHR_0_io_mem_req_bits_client_xact_id ),
       //.io_in_0_bits_data(  )
       .io_in_0_bits_a_type( MSHR_0_io_mem_req_bits_a_type ),
       //.io_in_0_bits_write_mask(  )
       //.io_in_0_bits_subword_addr(  )
       //.io_in_0_bits_atomic_opcode(  )
       .io_out_ready( io_mem_req_ready ),
       .io_out_valid( mem_req_arb_io_out_valid ),
       .io_out_bits_addr( mem_req_arb_io_out_bits_addr ),
       .io_out_bits_client_xact_id( mem_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_data( mem_req_arb_io_out_bits_data ),
       .io_out_bits_a_type( mem_req_arb_io_out_bits_a_type ),
       .io_out_bits_write_mask( mem_req_arb_io_out_bits_write_mask ),
       .io_out_bits_subword_addr( mem_req_arb_io_out_bits_subword_addr ),
       .io_out_bits_atomic_opcode( mem_req_arb_io_out_bits_atomic_opcode )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign mem_req_arb.io_in_1_bits_data = {16{$random}};
    assign mem_req_arb.io_in_1_bits_write_mask = {1{$random}};
    assign mem_req_arb.io_in_1_bits_subword_addr = {1{$random}};
    assign mem_req_arb.io_in_1_bits_atomic_opcode = {1{$random}};
    assign mem_req_arb.io_in_0_bits_data = {16{$random}};
    assign mem_req_arb.io_in_0_bits_write_mask = {1{$random}};
    assign mem_req_arb.io_in_0_bits_subword_addr = {1{$random}};
    assign mem_req_arb.io_in_0_bits_atomic_opcode = {1{$random}};
  `endif
  Arbiter_3 mem_finish_arb(
       .io_in_1_ready( mem_finish_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_finish_valid ),
       .io_in_1_bits_header_src( MSHR_1_io_mem_finish_bits_header_src ),
       .io_in_1_bits_header_dst( MSHR_1_io_mem_finish_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( MSHR_1_io_mem_finish_bits_payload_master_xact_id ),
       .io_in_0_ready( mem_finish_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_mem_finish_valid ),
       .io_in_0_bits_header_src( MSHR_0_io_mem_finish_bits_header_src ),
       .io_in_0_bits_header_dst( MSHR_0_io_mem_finish_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( MSHR_0_io_mem_finish_bits_payload_master_xact_id ),
       .io_out_ready( io_mem_finish_ready ),
       .io_out_valid( mem_finish_arb_io_out_valid ),
       .io_out_bits_header_src( mem_finish_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( mem_finish_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( mem_finish_arb_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
  Arbiter_4 wb_req_arb(
       .io_in_1_ready( wb_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_wb_req_valid ),
       .io_in_1_bits_tag( MSHR_1_io_wb_req_bits_tag ),
       .io_in_1_bits_idx( MSHR_1_io_wb_req_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_master_xact_id( MSHR_1_io_wb_req_bits_master_xact_id ),
       .io_in_1_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_in_0_ready( wb_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_wb_req_valid ),
       .io_in_0_bits_tag( MSHR_0_io_wb_req_bits_tag ),
       .io_in_0_bits_idx( MSHR_0_io_wb_req_bits_idx ),
       .io_in_0_bits_way_en( MSHR_0_io_wb_req_bits_way_en ),
       .io_in_0_bits_client_xact_id( MSHR_0_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_master_xact_id( MSHR_0_io_wb_req_bits_master_xact_id ),
       .io_in_0_bits_r_type( MSHR_0_io_wb_req_bits_r_type ),
       .io_out_ready( io_wb_req_ready ),
       .io_out_valid( wb_req_arb_io_out_valid ),
       .io_out_bits_tag( wb_req_arb_io_out_bits_tag ),
       .io_out_bits_idx( wb_req_arb_io_out_bits_idx ),
       .io_out_bits_way_en( wb_req_arb_io_out_bits_way_en ),
       .io_out_bits_client_xact_id( wb_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_master_xact_id( wb_req_arb_io_out_bits_master_xact_id ),
       .io_out_bits_r_type( wb_req_arb_io_out_bits_r_type )
       //.io_chosen(  )
  );
  Arbiter_5 replay_arb(
       .io_in_1_ready( replay_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_replay_valid ),
       .io_in_1_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_in_1_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_in_1_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_in_1_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_in_1_bits_data( MSHR_1_io_replay_bits_data ),
       .io_in_1_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_in_1_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_in_1_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_in_0_ready( replay_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_replay_valid ),
       .io_in_0_bits_kill( MSHR_0_io_replay_bits_kill ),
       .io_in_0_bits_typ( MSHR_0_io_replay_bits_typ ),
       .io_in_0_bits_phys( MSHR_0_io_replay_bits_phys ),
       .io_in_0_bits_addr( MSHR_0_io_replay_bits_addr ),
       .io_in_0_bits_data( MSHR_0_io_replay_bits_data ),
       .io_in_0_bits_tag( MSHR_0_io_replay_bits_tag ),
       .io_in_0_bits_cmd( MSHR_0_io_replay_bits_cmd ),
       .io_in_0_bits_sdq_id( MSHR_0_io_replay_bits_sdq_id ),
       .io_out_ready( io_replay_ready ),
       .io_out_valid( replay_arb_io_out_valid ),
       .io_out_bits_kill( replay_arb_io_out_bits_kill ),
       .io_out_bits_typ( replay_arb_io_out_bits_typ ),
       .io_out_bits_phys( replay_arb_io_out_bits_phys ),
       .io_out_bits_addr( replay_arb_io_out_bits_addr ),
       //.io_out_bits_data(  )
       .io_out_bits_tag( replay_arb_io_out_bits_tag ),
       .io_out_bits_cmd( replay_arb_io_out_bits_cmd ),
       .io_out_bits_sdq_id( replay_arb_io_out_bits_sdq_id )
       //.io_chosen(  )
  );
  Arbiter_6 alloc_arb(
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_req_pri_rdy ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_req_pri_rdy ),
       //.io_in_0_bits(  )
       .io_out_ready( T114 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
  `endif
  MSHR_0 MSHR_0(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_0_ready ),
       .io_req_pri_rdy( MSHR_0_io_req_pri_rdy ),
       .io_req_sec_val( T112 ),
       .io_req_sec_rdy( MSHR_0_io_req_sec_rdy ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_data( io_req_bits_data ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_req_sdq_id( T0 ),
       .io_idx_match( MSHR_0_io_idx_match ),
       .io_tag( MSHR_0_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_0_ready ),
       .io_mem_req_valid( MSHR_0_io_mem_req_valid ),
       .io_mem_req_bits_addr( MSHR_0_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( MSHR_0_io_mem_req_bits_client_xact_id ),
       //.io_mem_req_bits_data(  )
       .io_mem_req_bits_a_type( MSHR_0_io_mem_req_bits_a_type ),
       //.io_mem_req_bits_write_mask(  )
       //.io_mem_req_bits_subword_addr(  )
       //.io_mem_req_bits_atomic_opcode(  )
       .io_mem_resp_way_en( MSHR_0_io_mem_resp_way_en ),
       .io_mem_resp_addr( MSHR_0_io_mem_resp_addr ),
       .io_mem_resp_wmask( MSHR_0_io_mem_resp_wmask ),
       .io_mem_resp_data( MSHR_0_io_mem_resp_data ),
       .io_meta_read_ready( meta_read_arb_io_in_0_ready ),
       .io_meta_read_valid( MSHR_0_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_0_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_0_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_0_ready ),
       .io_meta_write_valid( MSHR_0_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_0_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_0_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_0_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_0_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_0_ready ),
       .io_replay_valid( MSHR_0_io_replay_valid ),
       .io_replay_bits_kill( MSHR_0_io_replay_bits_kill ),
       .io_replay_bits_typ( MSHR_0_io_replay_bits_typ ),
       .io_replay_bits_phys( MSHR_0_io_replay_bits_phys ),
       .io_replay_bits_addr( MSHR_0_io_replay_bits_addr ),
       .io_replay_bits_data( MSHR_0_io_replay_bits_data ),
       .io_replay_bits_tag( MSHR_0_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_0_io_replay_bits_cmd ),
       .io_replay_bits_sdq_id( MSHR_0_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( mem_finish_arb_io_in_0_ready ),
       .io_mem_finish_valid( MSHR_0_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( MSHR_0_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( MSHR_0_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( MSHR_0_io_mem_finish_bits_payload_master_xact_id ),
       .io_wb_req_ready( wb_req_arb_io_in_0_ready ),
       .io_wb_req_valid( MSHR_0_io_wb_req_valid ),
       .io_wb_req_bits_tag( MSHR_0_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( MSHR_0_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( MSHR_0_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( MSHR_0_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( MSHR_0_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( MSHR_0_io_wb_req_bits_r_type ),
       .io_probe_rdy( MSHR_0_io_probe_rdy )
  );
  `ifndef SYNTHESIS
    assign MSHR_0.io_mem_resp_wmask = {1{$random}};
  `endif
  MSHR_1 MSHR_1(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_1_ready ),
       .io_req_pri_rdy( MSHR_1_io_req_pri_rdy ),
       .io_req_sec_val( T104 ),
       .io_req_sec_rdy( MSHR_1_io_req_sec_rdy ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_data( io_req_bits_data ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_req_sdq_id( T0 ),
       .io_idx_match( MSHR_1_io_idx_match ),
       .io_tag( MSHR_1_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_1_ready ),
       .io_mem_req_valid( MSHR_1_io_mem_req_valid ),
       .io_mem_req_bits_addr( MSHR_1_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       //.io_mem_req_bits_data(  )
       .io_mem_req_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       //.io_mem_req_bits_write_mask(  )
       //.io_mem_req_bits_subword_addr(  )
       //.io_mem_req_bits_atomic_opcode(  )
       .io_mem_resp_way_en( MSHR_1_io_mem_resp_way_en ),
       .io_mem_resp_addr( MSHR_1_io_mem_resp_addr ),
       .io_mem_resp_wmask( MSHR_1_io_mem_resp_wmask ),
       .io_mem_resp_data( MSHR_1_io_mem_resp_data ),
       .io_meta_read_ready( meta_read_arb_io_in_1_ready ),
       .io_meta_read_valid( MSHR_1_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_1_ready ),
       .io_meta_write_valid( MSHR_1_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_1_ready ),
       .io_replay_valid( MSHR_1_io_replay_valid ),
       .io_replay_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_replay_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_replay_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_replay_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_replay_bits_data( MSHR_1_io_replay_bits_data ),
       .io_replay_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_replay_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( mem_finish_arb_io_in_1_ready ),
       .io_mem_finish_valid( MSHR_1_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( MSHR_1_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( MSHR_1_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( MSHR_1_io_mem_finish_bits_payload_master_xact_id ),
       .io_wb_req_ready( wb_req_arb_io_in_1_ready ),
       .io_wb_req_valid( MSHR_1_io_wb_req_valid ),
       .io_wb_req_bits_tag( MSHR_1_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( MSHR_1_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( MSHR_1_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_probe_rdy( MSHR_1_io_probe_rdy )
  );
  `ifndef SYNTHESIS
    assign MSHR_1.io_mem_resp_wmask = {1{$random}};
  `endif

  always @(posedge clk) begin
    sdq_val <= T19;
    if(free_sdq) begin
      R130 <= replay_arb_io_out_bits_sdq_id;
    end
  end
endmodule

module MetadataArray(input clk, input reset,
    output io_read_ready,
    input  io_read_valid,
    input [5:0] io_read_bits_idx,
    output io_write_ready,
    input  io_write_valid,
    input [5:0] io_write_bits_idx,
    input  io_write_bits_way_en,
    input [19:0] io_write_bits_data_tag,
    input [1:0] io_write_bits_data_coh_state,
    output[19:0] io_resp_0_tag,
    output[1:0] io_resp_0_coh_state
);

  wire[1:0] T0;
  wire[21:0] T1;
  wire[21:0] T2;
  reg [21:0] tag_arr [63:0];
  wire[21:0] T3;
  wire[21:0] T4;
  wire[21:0] T5;
  wire[21:0] T6;
  wire[21:0] T7;
  wire[21:0] T8;
  wire[21:0] T9;
  wire T10;
  wire wmask;
  wire T11;
  reg [6:0] rst_cnt;
  wire[6:0] T12;
  wire[6:0] T13;
  wire[6:0] T14;
  wire[21:0] T15;
  wire[5:0] T16;
  wire[6:0] waddr;
  wire[6:0] T17;
  wire[21:0] T18;
  wire[21:0] wdata;
  wire[21:0] T19;
  wire[1:0] T20;
  wire[21:0] T21;
  wire[21:0] T22;
  wire[21:0] T23;
  wire[1:0] rstVal_coh_state;
  wire[1:0] T24;
  wire[19:0] rstVal_tag;
  wire[19:0] T25;
  wire T26;
  wire[5:0] T27;
  reg [5:0] R28;
  wire[5:0] T29;
  wire[19:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 64; initvar = initvar+1)
      tag_arr[initvar] = {1{$random}};
    rst_cnt = {1{$random}};
    R28 = {1{$random}};
  end
`endif

  assign io_resp_0_coh_state = T0;
  assign T0 = T1[1'h1:1'h0];
  assign T1 = T2[5'h15:1'h0];
  assign T2 = tag_arr[R28];
  always @(posedge clk)
    if (T26)
      tag_arr[T27] <= T4;
  assign T4 = T18 | T5;
  assign T5 = T15 & T6;
  assign T6 = ~ T7;
  assign T7 = T8;
  assign T8 = 22'h0 - T9;
  assign T9 = {21'h0, T10};
  assign T10 = wmask;
  assign wmask = T11 ? 1'h1 : io_write_bits_way_en;
  assign T11 = rst_cnt < 7'h40;
  assign T12 = reset ? 7'h0 : T13;
  assign T13 = T11 ? T14 : rst_cnt;
  assign T14 = rst_cnt + 7'h1;
  assign T15 = tag_arr[T16];
  assign T16 = waddr[3'h5:1'h0];
  assign waddr = T11 ? rst_cnt : T17;
  assign T17 = {1'h0, io_write_bits_idx};
  assign T18 = wdata & T7;
  assign wdata = T19;
  assign T19 = {T25, T20};
  assign T20 = T21[1'h1:1'h0];
  assign T21 = T11 ? T23 : T22;
  assign T22 = {io_write_bits_data_tag, io_write_bits_data_coh_state};
  assign T23 = {rstVal_tag, rstVal_coh_state};
  assign rstVal_coh_state = T24;
  assign T24 = 2'h0;
  assign rstVal_tag = 20'h0;
  assign T25 = T21[5'h15:2'h2];
  assign T26 = T11 | io_write_valid;
  assign T27 = waddr[3'h5:1'h0];
  assign T29 = io_read_valid ? io_read_bits_idx : R28;
  assign io_resp_0_tag = T30;
  assign T30 = T1[5'h15:2'h2];
  assign io_write_ready = T31;
  assign T31 = T11 ^ 1'h1;
  assign io_read_ready = T32;
  assign T32 = T34 & T33;
  assign T33 = io_write_valid ^ 1'h1;
  assign T34 = T11 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      rst_cnt <= 7'h0;
    end else if(T11) begin
      rst_cnt <= T14;
    end
    if(io_read_valid) begin
      R28 <= io_read_bits_idx;
    end
  end
endmodule

module Arbiter_7(
    output io_in_4_ready,
    input  io_in_4_valid,
    input [5:0] io_in_4_bits_idx,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [5:0] io_in_3_bits_idx,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [5:0] io_in_2_bits_idx,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[5:0] T5;
  wire[5:0] T6;
  wire[5:0] T7;
  wire T8;
  wire[2:0] T9;
  wire[5:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : 3'h4;
  assign io_out_bits_idx = T5;
  assign T5 = T13 ? io_in_4_bits_idx : T6;
  assign T6 = T12 ? T10 : T7;
  assign T7 = T8 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign T8 = T9[1'h0:1'h0];
  assign T9 = T0;
  assign T10 = T11 ? io_in_3_bits_idx : io_in_2_bits_idx;
  assign T11 = T9[1'h0:1'h0];
  assign T12 = T9[1'h1:1'h1];
  assign T13 = T9[2'h2:2'h2];
  assign io_out_valid = T14;
  assign T14 = T21 ? io_in_4_valid : T15;
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? io_in_1_valid : io_in_0_valid;
  assign T17 = T9[1'h0:1'h0];
  assign T18 = T19 ? io_in_3_valid : io_in_2_valid;
  assign T19 = T9[1'h0:1'h0];
  assign T20 = T9[1'h1:1'h1];
  assign T21 = T9[2'h2:2'h2];
  assign io_in_0_ready = T22;
  assign T22 = T23 & io_out_ready;
  assign T23 = 1'h1;
  assign io_in_1_ready = T24;
  assign T24 = T25 & io_out_ready;
  assign T25 = T26;
  assign T26 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T27;
  assign T27 = T28 & io_out_ready;
  assign T28 = T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T31;
  assign T31 = T32 & io_out_ready;
  assign T32 = T33;
  assign T33 = T34 ^ 1'h1;
  assign T34 = T35 | io_in_2_valid;
  assign T35 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T36;
  assign T36 = T37 & io_out_ready;
  assign T37 = T38;
  assign T38 = T39 ^ 1'h1;
  assign T39 = T40 | io_in_3_valid;
  assign T40 = T41 | io_in_2_valid;
  assign T41 = io_in_0_valid | io_in_1_valid;
endmodule

module DataArray(input clk,
    output io_read_ready,
    input  io_read_valid,
    input  io_read_bits_way_en,
    input [11:0] io_read_bits_addr,
    output io_write_ready,
    input  io_write_valid,
    input  io_write_bits_way_en,
    input [11:0] io_write_bits_addr,
    input [1:0] io_write_bits_wmask,
    input [127:0] io_write_bits_data,
    output[127:0] io_resp_0
);

  wire[127:0] T0;
  reg [127:0] T1 [255:0];
  wire[127:0] T2;
  wire[127:0] T3;
  wire[127:0] T4;
  wire[127:0] T5;
  wire[127:0] T6;
  wire[127:0] T7;
  wire[63:0] T8;
  wire[63:0] T9;
  wire T10;
  wire[63:0] T11;
  wire[63:0] T12;
  wire T13;
  wire[127:0] T14;
  wire[7:0] waddr;
  wire[127:0] T15;
  wire T16;
  reg [7:0] R17;
  wire[7:0] T18;
  wire[7:0] raddr;
  wire T19;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 256; initvar = initvar+1)
      T1[initvar] = {4{$random}};
    R17 = {1{$random}};
  end
`endif

  assign io_resp_0 = T0;
  assign T0 = T1[R17];
  always @(posedge clk)
    if (T16)
      T1[waddr] <= T3;
  assign T3 = T15 | T4;
  assign T4 = T14 & T5;
  assign T5 = ~ T6;
  assign T6 = T7;
  assign T7 = {T11, T8};
  assign T8 = 64'h0 - T9;
  assign T9 = {63'h0, T10};
  assign T10 = io_write_bits_wmask[1'h0:1'h0];
  assign T11 = 64'h0 - T12;
  assign T12 = {63'h0, T13};
  assign T13 = io_write_bits_wmask[1'h1:1'h1];
  assign T14 = T1[waddr];
  assign waddr = io_write_bits_addr >> 3'h4;
  assign T15 = io_write_bits_data & T6;
  assign T16 = io_write_bits_way_en & io_write_valid;
  assign T18 = T19 ? raddr : R17;
  assign raddr = io_read_bits_addr >> 3'h4;
  assign T19 = io_read_bits_way_en & io_read_valid;
  assign io_write_ready = 1'h1;
  assign io_read_ready = 1'h1;

  always @(posedge clk) begin
    if(T19) begin
      R17 <= raddr;
    end
  end
endmodule

module Arbiter_8(
    output io_in_3_ready,
    input  io_in_3_valid,
    input  io_in_3_bits_way_en,
    input [11:0] io_in_3_bits_addr,
    output io_in_2_ready,
    input  io_in_2_valid,
    input  io_in_2_bits_way_en,
    input [11:0] io_in_2_bits_addr,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_way_en,
    input [11:0] io_in_1_bits_addr,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_way_en,
    input [11:0] io_in_0_bits_addr,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_way_en,
    output[11:0] io_out_bits_addr,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[11:0] T4;
  wire[11:0] T5;
  wire T6;
  wire[1:0] T7;
  wire[11:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 2'h0 : T2;
  assign T2 = io_in_1_valid ? 2'h1 : T3;
  assign T3 = io_in_2_valid ? 2'h2 : 2'h3;
  assign io_out_bits_addr = T4;
  assign T4 = T10 ? T8 : T5;
  assign T5 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign T6 = T7[1'h0:1'h0];
  assign T7 = T0;
  assign T8 = T9 ? io_in_3_bits_addr : io_in_2_bits_addr;
  assign T9 = T7[1'h0:1'h0];
  assign T10 = T7[1'h1:1'h1];
  assign io_out_bits_way_en = T11;
  assign T11 = T16 ? T14 : T12;
  assign T12 = T13 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign T13 = T7[1'h0:1'h0];
  assign T14 = T15 ? io_in_3_bits_way_en : io_in_2_bits_way_en;
  assign T15 = T7[1'h0:1'h0];
  assign T16 = T7[1'h1:1'h1];
  assign io_out_valid = T17;
  assign T17 = T22 ? T20 : T18;
  assign T18 = T19 ? io_in_1_valid : io_in_0_valid;
  assign T19 = T7[1'h0:1'h0];
  assign T20 = T21 ? io_in_3_valid : io_in_2_valid;
  assign T21 = T7[1'h0:1'h0];
  assign T22 = T7[1'h1:1'h1];
  assign io_in_0_ready = T23;
  assign T23 = T24 & io_out_ready;
  assign T24 = 1'h1;
  assign io_in_1_ready = T25;
  assign T25 = T26 & io_out_ready;
  assign T26 = T27;
  assign T27 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T28;
  assign T28 = T29 & io_out_ready;
  assign T29 = T30;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T32;
  assign T32 = T33 & io_out_ready;
  assign T33 = T34;
  assign T34 = T35 ^ 1'h1;
  assign T35 = T36 | io_in_2_valid;
  assign T36 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_9(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_way_en,
    input [11:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_wmask,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_way_en,
    input [11:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_wmask,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_way_en,
    output[11:0] io_out_bits_addr,
    output[1:0] io_out_bits_wmask,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[127:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[11:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_data = T2;
  assign T2 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T3 = T0;
  assign io_out_bits_wmask = T4;
  assign T4 = T3 ? io_in_1_bits_wmask : io_in_0_bits_wmask;
  assign io_out_bits_addr = T5;
  assign T5 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_way_en = T6;
  assign T6 = T3 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_valid = T7;
  assign T7 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T8;
  assign T8 = T9 & io_out_ready;
  assign T9 = 1'h1;
  assign io_in_1_ready = T10;
  assign T10 = T11 & io_out_ready;
  assign T11 = T12;
  assign T12 = io_in_0_valid ^ 1'h1;
endmodule

module AMOALU(
    input [5:0] io_addr,
    input [3:0] io_cmd,
    input [2:0] io_typ,
    input [63:0] io_lhs,
    input [63:0] io_rhs,
    output[63:0] io_out
);

  wire[63:0] T0;
  wire[87:0] T1;
  wire[87:0] T2;
  wire[87:0] T3;
  wire[87:0] T4;
  wire[87:0] wmask;
  wire[87:0] T5;
  wire[47:0] T6;
  wire[23:0] T7;
  wire[15:0] T8;
  wire[7:0] T9;
  wire[7:0] T10;
  wire T11;
  wire[10:0] T12;
  wire[10:0] T13;
  wire[10:0] T14;
  wire[10:0] T15;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[10:0] T21;
  wire[8:0] T22;
  wire[2:0] T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire T27;
  wire[10:0] T28;
  wire[7:0] T29;
  wire[2:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire[7:0] T35;
  wire T36;
  wire[7:0] T37;
  wire[7:0] T38;
  wire T39;
  wire[23:0] T40;
  wire[15:0] T41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire T44;
  wire[7:0] T45;
  wire[7:0] T46;
  wire T47;
  wire[7:0] T48;
  wire[7:0] T49;
  wire T50;
  wire[39:0] T51;
  wire[23:0] T52;
  wire[15:0] T53;
  wire[7:0] T54;
  wire[7:0] T55;
  wire T56;
  wire[7:0] T57;
  wire[7:0] T58;
  wire T59;
  wire[7:0] T60;
  wire[7:0] T61;
  wire T62;
  wire[15:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire T69;
  wire[87:0] T70;
  wire[87:0] T71;
  wire[63:0] out;
  wire[63:0] T72;
  wire[63:0] T73;
  wire[63:0] T74;
  wire[63:0] T75;
  wire[63:0] T76;
  wire[63:0] T77;
  wire[63:0] rhs;
  wire[63:0] T78;
  wire[31:0] T79;
  wire[63:0] T80;
  wire[31:0] T81;
  wire[15:0] T82;
  wire[63:0] T83;
  wire[31:0] T84;
  wire[15:0] T85;
  wire[7:0] T86;
  wire T87;
  wire max;
  wire T88;
  wire[4:0] T89;
  wire T90;
  wire[4:0] T91;
  wire min;
  wire T92;
  wire[4:0] T93;
  wire T94;
  wire[4:0] T95;
  wire less;
  wire T96;
  wire cmp_rhs;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire word;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire cmp_lhs;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire sgned;
  wire T113;
  wire[4:0] T114;
  wire T115;
  wire[4:0] T116;
  wire lt;
  wire T117;
  wire T118;
  wire T119;
  wire[31:0] T120;
  wire[31:0] T121;
  wire eq_hi;
  wire[31:0] T122;
  wire[31:0] T123;
  wire T124;
  wire[31:0] T125;
  wire[31:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire[63:0] T130;
  wire T131;
  wire[4:0] T132;
  wire[63:0] T133;
  wire T134;
  wire[4:0] T135;
  wire[63:0] T136;
  wire T137;
  wire[4:0] T138;
  wire[63:0] adder_out;
  wire[63:0] T139;
  wire[63:0] mask;
  wire[63:0] T140;
  wire[31:0] T141;
  wire T142;
  wire[63:0] T143;
  wire[63:0] T144;
  wire T145;
  wire[4:0] T146;


  assign io_out = T0;
  assign T0 = T1[6'h3f:1'h0];
  assign T1 = T70 | T2;
  assign T2 = T4 & T3;
  assign T3 = {24'h0, io_lhs};
  assign T4 = ~ wmask;
  assign wmask = T5;
  assign T5 = {T51, T6};
  assign T6 = {T40, T7};
  assign T7 = {T37, T8};
  assign T8 = {T34, T9};
  assign T9 = 8'h0 - T10;
  assign T10 = {7'h0, T11};
  assign T11 = T12[1'h0:1'h0];
  assign T12 = T31 ? T28 : T13;
  assign T13 = T25 ? T21 : T14;
  assign T14 = T18 ? T15 : 11'hff;
  assign T15 = 4'hf << T16;
  assign T16 = {T17, 2'h0};
  assign T17 = io_addr[2'h2:2'h2];
  assign T18 = T20 | T19;
  assign T19 = io_typ == 3'h6;
  assign T20 = io_typ == 3'h2;
  assign T21 = {2'h0, T22};
  assign T22 = 2'h3 << T23;
  assign T23 = {T24, 1'h0};
  assign T24 = io_addr[2'h2:1'h1];
  assign T25 = T27 | T26;
  assign T26 = io_typ == 3'h5;
  assign T27 = io_typ == 3'h1;
  assign T28 = {3'h0, T29};
  assign T29 = 1'h1 << T30;
  assign T30 = io_addr[2'h2:1'h0];
  assign T31 = T33 | T32;
  assign T32 = io_typ == 3'h4;
  assign T33 = io_typ == 3'h0;
  assign T34 = 8'h0 - T35;
  assign T35 = {7'h0, T36};
  assign T36 = T12[1'h1:1'h1];
  assign T37 = 8'h0 - T38;
  assign T38 = {7'h0, T39};
  assign T39 = T12[2'h2:2'h2];
  assign T40 = {T48, T41};
  assign T41 = {T45, T42};
  assign T42 = 8'h0 - T43;
  assign T43 = {7'h0, T44};
  assign T44 = T12[2'h3:2'h3];
  assign T45 = 8'h0 - T46;
  assign T46 = {7'h0, T47};
  assign T47 = T12[3'h4:3'h4];
  assign T48 = 8'h0 - T49;
  assign T49 = {7'h0, T50};
  assign T50 = T12[3'h5:3'h5];
  assign T51 = {T63, T52};
  assign T52 = {T60, T53};
  assign T53 = {T57, T54};
  assign T54 = 8'h0 - T55;
  assign T55 = {7'h0, T56};
  assign T56 = T12[3'h6:3'h6];
  assign T57 = 8'h0 - T58;
  assign T58 = {7'h0, T59};
  assign T59 = T12[3'h7:3'h7];
  assign T60 = 8'h0 - T61;
  assign T61 = {7'h0, T62};
  assign T62 = T12[4'h8:4'h8];
  assign T63 = {T67, T64};
  assign T64 = 8'h0 - T65;
  assign T65 = {7'h0, T66};
  assign T66 = T12[4'h9:4'h9];
  assign T67 = 8'h0 - T68;
  assign T68 = {7'h0, T69};
  assign T69 = T12[4'ha:4'ha];
  assign T70 = wmask & T71;
  assign T71 = {24'h0, out};
  assign out = T145 ? adder_out : T72;
  assign T72 = T137 ? T136 : T73;
  assign T73 = T134 ? T133 : T74;
  assign T74 = T131 ? T130 : T75;
  assign T75 = T87 ? io_lhs : T76;
  assign T76 = T31 ? T83 : T77;
  assign T77 = T25 ? T80 : rhs;
  assign rhs = T18 ? T78 : io_rhs;
  assign T78 = {T79, T79};
  assign T79 = io_rhs[5'h1f:1'h0];
  assign T80 = {T81, T81};
  assign T81 = {T82, T82};
  assign T82 = io_rhs[4'hf:1'h0];
  assign T83 = {T84, T84};
  assign T84 = {T85, T85};
  assign T85 = {T86, T86};
  assign T86 = io_rhs[3'h7:1'h0];
  assign T87 = less ? min : max;
  assign max = T90 | T88;
  assign T88 = T89 == 5'hf;
  assign T89 = {1'h0, io_cmd};
  assign T90 = T91 == 5'hd;
  assign T91 = {1'h0, io_cmd};
  assign min = T94 | T92;
  assign T92 = T93 == 5'he;
  assign T93 = {1'h0, io_cmd};
  assign T94 = T95 == 5'hc;
  assign T95 = {1'h0, io_cmd};
  assign less = T129 ? lt : T96;
  assign T96 = sgned ? cmp_lhs : cmp_rhs;
  assign cmp_rhs = T99 ? T98 : T97;
  assign T97 = rhs[6'h3f:6'h3f];
  assign T98 = rhs[5'h1f:5'h1f];
  assign T99 = word & T100;
  assign T100 = T101 ^ 1'h1;
  assign T101 = io_addr[2'h2:2'h2];
  assign word = T103 | T102;
  assign T102 = io_typ == 3'h4;
  assign T103 = T105 | T104;
  assign T104 = io_typ == 3'h0;
  assign T105 = T107 | T106;
  assign T106 = io_typ == 3'h6;
  assign T107 = io_typ == 3'h2;
  assign cmp_lhs = T110 ? T109 : T108;
  assign T108 = io_lhs[6'h3f:6'h3f];
  assign T109 = io_lhs[5'h1f:5'h1f];
  assign T110 = word & T111;
  assign T111 = T112 ^ 1'h1;
  assign T112 = io_addr[2'h2:2'h2];
  assign sgned = T115 | T113;
  assign T113 = T114 == 5'hd;
  assign T114 = {1'h0, io_cmd};
  assign T115 = T116 == 5'hc;
  assign T116 = {1'h0, io_cmd};
  assign lt = word ? T127 : T117;
  assign T117 = T124 | T118;
  assign T118 = eq_hi & T119;
  assign T119 = T121 < T120;
  assign T120 = rhs[5'h1f:1'h0];
  assign T121 = io_lhs[5'h1f:1'h0];
  assign eq_hi = T123 == T122;
  assign T122 = rhs[6'h3f:6'h20];
  assign T123 = io_lhs[6'h3f:6'h20];
  assign T124 = T126 < T125;
  assign T125 = rhs[6'h3f:6'h20];
  assign T126 = io_lhs[6'h3f:6'h20];
  assign T127 = T128 ? T124 : T119;
  assign T128 = io_addr[2'h2:2'h2];
  assign T129 = cmp_lhs == cmp_rhs;
  assign T130 = io_lhs ^ rhs;
  assign T131 = T132 == 5'h9;
  assign T132 = {1'h0, io_cmd};
  assign T133 = io_lhs | rhs;
  assign T134 = T135 == 5'ha;
  assign T135 = {1'h0, io_cmd};
  assign T136 = io_lhs & rhs;
  assign T137 = T138 == 5'hb;
  assign T138 = {1'h0, io_cmd};
  assign adder_out = T143 + T139;
  assign T139 = rhs & mask;
  assign mask = 64'hffffffffffffffff ^ T140;
  assign T140 = {32'h0, T141};
  assign T141 = T142 << 5'h1f;
  assign T142 = io_addr[2'h2:2'h2];
  assign T143 = T144;
  assign T144 = io_lhs & mask;
  assign T145 = T146 == 5'h8;
  assign T146 = {1'h0, io_cmd};
endmodule

module Arbiter_10(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr,
    input [3:0] io_in_1_bits_client_xact_id,
    input [3:0] io_in_1_bits_master_xact_id,
    input [511:0] io_in_1_bits_data,
    input [2:0] io_in_1_bits_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr,
    input [3:0] io_in_0_bits_client_xact_id,
    input [3:0] io_in_0_bits_master_xact_id,
    input [511:0] io_in_0_bits_data,
    input [2:0] io_in_0_bits_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr,
    output[3:0] io_out_bits_client_xact_id,
    output[3:0] io_out_bits_master_xact_id,
    output[511:0] io_out_bits_data,
    output[2:0] io_out_bits_r_type,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[2:0] T2;
  wire T3;
  wire[511:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[25:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_r_type = T2;
  assign T2 = T3 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign T3 = T0;
  assign io_out_bits_data = T4;
  assign T4 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_master_xact_id = T5;
  assign T5 = T3 ? io_in_1_bits_master_xact_id : io_in_0_bits_master_xact_id;
  assign io_out_bits_client_xact_id = T6;
  assign T6 = T3 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr = T7;
  assign T7 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T8;
  assign T8 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = 1'h1;
  assign io_in_1_ready = T11;
  assign T11 = T12 & io_out_ready;
  assign T12 = T13;
  assign T13 = io_in_0_valid ^ 1'h1;
endmodule

module FlowThroughSerializer_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [1:0] io_in_bits_header_src,
    input [1:0] io_in_bits_header_dst,
    input [511:0] io_in_bits_payload_data,
    input [3:0] io_in_bits_payload_client_xact_id,
    input [3:0] io_in_bits_payload_master_xact_id,
    input [3:0] io_in_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[3:0] io_out_bits_payload_client_xact_id,
    output[3:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[1:0] io_cnt,
    output io_done
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg  active;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire wrap;
  reg [1:0] cnt;
  wire[1:0] T16;
  wire[1:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire[3:0] T23;
  reg [3:0] rbits_payload_g_type;
  wire[3:0] T24;
  wire[3:0] T25;
  wire[3:0] T26;
  reg [3:0] rbits_payload_master_xact_id;
  wire[3:0] T27;
  wire[3:0] T28;
  wire[3:0] T29;
  reg [3:0] rbits_payload_client_xact_id;
  wire[3:0] T30;
  wire[3:0] T31;
  wire[511:0] T32;
  wire[511:0] T33;
  reg [511:0] rbits_payload_data;
  wire[511:0] T34;
  wire[511:0] T35;
  wire[511:0] T36;
  wire[127:0] T37;
  wire[127:0] T38;
  wire[127:0] shifter_0;
  wire[127:0] T39;
  wire[127:0] shifter_1;
  wire[127:0] T40;
  wire T41;
  wire[1:0] T42;
  wire[127:0] T43;
  wire[127:0] shifter_2;
  wire[127:0] T44;
  wire[127:0] shifter_3;
  wire[127:0] T45;
  wire T46;
  wire T47;
  wire[1:0] T48;
  reg [1:0] rbits_header_dst;
  wire[1:0] T49;
  wire[1:0] T50;
  wire[1:0] T51;
  reg [1:0] rbits_header_src;
  wire[1:0] T52;
  wire[1:0] T53;
  wire T54;
  wire T55;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    active = {1{$random}};
    cnt = {1{$random}};
    rbits_payload_g_type = {1{$random}};
    rbits_payload_master_xact_id = {1{$random}};
    rbits_payload_client_xact_id = {1{$random}};
    rbits_payload_data = {16{$random}};
    rbits_header_dst = {1{$random}};
    rbits_header_src = {1{$random}};
  end
`endif

  assign io_done = T0;
  assign T0 = T15 ? 1'h1 : T1;
  assign T1 = T6 ? T2 : 1'h0;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 | T4;
  assign T4 = io_in_bits_payload_g_type == 4'h2;
  assign T5 = io_in_bits_payload_g_type == 4'h1;
  assign T6 = T7 & io_in_valid;
  assign T7 = active ^ 1'h1;
  assign T8 = reset ? 1'h0 : T9;
  assign T9 = T15 ? 1'h0 : T10;
  assign T10 = T11 ? 1'h1 : active;
  assign T11 = T6 & T12;
  assign T12 = T14 | T13;
  assign T13 = io_in_bits_payload_g_type == 4'h2;
  assign T14 = io_in_bits_payload_g_type == 4'h1;
  assign T15 = T22 & wrap;
  assign wrap = cnt == 2'h3;
  assign T16 = reset ? 2'h0 : T17;
  assign T17 = T15 ? 2'h0 : T18;
  assign T18 = T22 ? T21 : T19;
  assign T19 = T11 ? T20 : cnt;
  assign T20 = {1'h0, io_out_ready};
  assign T21 = cnt + 2'h1;
  assign T22 = active & io_out_ready;
  assign io_cnt = cnt;
  assign io_out_bits_payload_g_type = T23;
  assign T23 = active ? rbits_payload_g_type : io_in_bits_payload_g_type;
  assign T24 = reset ? io_in_bits_payload_g_type : T25;
  assign T25 = T11 ? io_in_bits_payload_g_type : rbits_payload_g_type;
  assign io_out_bits_payload_master_xact_id = T26;
  assign T26 = active ? rbits_payload_master_xact_id : io_in_bits_payload_master_xact_id;
  assign T27 = reset ? io_in_bits_payload_master_xact_id : T28;
  assign T28 = T11 ? io_in_bits_payload_master_xact_id : rbits_payload_master_xact_id;
  assign io_out_bits_payload_client_xact_id = T29;
  assign T29 = active ? rbits_payload_client_xact_id : io_in_bits_payload_client_xact_id;
  assign T30 = reset ? io_in_bits_payload_client_xact_id : T31;
  assign T31 = T11 ? io_in_bits_payload_client_xact_id : rbits_payload_client_xact_id;
  assign io_out_bits_payload_data = T32;
  assign T32 = active ? T36 : T33;
  assign T33 = active ? rbits_payload_data : io_in_bits_payload_data;
  assign T34 = reset ? io_in_bits_payload_data : T35;
  assign T35 = T11 ? io_in_bits_payload_data : rbits_payload_data;
  assign T36 = {384'h0, T37};
  assign T37 = T47 ? T43 : T38;
  assign T38 = T41 ? shifter_1 : shifter_0;
  assign shifter_0 = T39;
  assign T39 = rbits_payload_data[7'h7f:1'h0];
  assign shifter_1 = T40;
  assign T40 = rbits_payload_data[8'hff:8'h80];
  assign T41 = T42[1'h0:1'h0];
  assign T42 = cnt;
  assign T43 = T46 ? shifter_3 : shifter_2;
  assign shifter_2 = T44;
  assign T44 = rbits_payload_data[9'h17f:9'h100];
  assign shifter_3 = T45;
  assign T45 = rbits_payload_data[9'h1ff:9'h180];
  assign T46 = T42[1'h0:1'h0];
  assign T47 = T42[1'h1:1'h1];
  assign io_out_bits_header_dst = T48;
  assign T48 = active ? rbits_header_dst : io_in_bits_header_dst;
  assign T49 = reset ? io_in_bits_header_dst : T50;
  assign T50 = T11 ? io_in_bits_header_dst : rbits_header_dst;
  assign io_out_bits_header_src = T51;
  assign T51 = active ? rbits_header_src : io_in_bits_header_src;
  assign T52 = reset ? io_in_bits_header_src : T53;
  assign T53 = T11 ? io_in_bits_header_src : rbits_header_src;
  assign io_out_valid = T54;
  assign T54 = active | io_in_valid;
  assign io_in_ready = T55;
  assign T55 = active ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      active <= 1'h0;
    end else if(T15) begin
      active <= 1'h0;
    end else if(T11) begin
      active <= 1'h1;
    end
    if(reset) begin
      cnt <= 2'h0;
    end else if(T15) begin
      cnt <= 2'h0;
    end else if(T22) begin
      cnt <= T21;
    end else if(T11) begin
      cnt <= T20;
    end
    if(reset) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end else if(T11) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end
    if(reset) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end else if(T11) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end
    if(reset) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end else if(T11) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end
    if(reset) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end else if(T11) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end
    if(reset) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end else if(T11) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end
    if(reset) begin
      rbits_header_src <= io_in_bits_header_src;
    end else if(T11) begin
      rbits_header_src <= io_in_bits_header_src;
    end
  end
endmodule

module HellaCache(input clk, input reset,
    output io_cpu_req_ready,
    input  io_cpu_req_valid,
    input  io_cpu_req_bits_kill,
    input [2:0] io_cpu_req_bits_typ,
    input  io_cpu_req_bits_phys,
    input [43:0] io_cpu_req_bits_addr,
    input [63:0] io_cpu_req_bits_data,
    input [7:0] io_cpu_req_bits_tag,
    input [4:0] io_cpu_req_bits_cmd,
    output io_cpu_resp_valid,
    output io_cpu_resp_bits_nack,
    output io_cpu_resp_bits_replay,
    output[2:0] io_cpu_resp_bits_typ,
    output io_cpu_resp_bits_has_data,
    output[63:0] io_cpu_resp_bits_data,
    output[63:0] io_cpu_resp_bits_data_subword,
    output[7:0] io_cpu_resp_bits_tag,
    output[3:0] io_cpu_resp_bits_cmd,
    output[43:0] io_cpu_resp_bits_addr,
    output[63:0] io_cpu_resp_bits_store_data,
    output io_cpu_replay_next_valid,
    output[7:0] io_cpu_replay_next_bits,
    output io_cpu_xcpt_ma_ld,
    output io_cpu_xcpt_ma_st,
    output io_cpu_xcpt_pf_ld,
    output io_cpu_xcpt_pf_st,
    input  io_cpu_ptw_req_ready,
    output io_cpu_ptw_req_valid,
    output[29:0] io_cpu_ptw_req_bits,
    input  io_cpu_ptw_resp_valid,
    input  io_cpu_ptw_resp_bits_error,
    input [18:0] io_cpu_ptw_resp_bits_ppn,
    input [5:0] io_cpu_ptw_resp_bits_perm,
    input [7:0] io_cpu_ptw_status_ip,
    input [7:0] io_cpu_ptw_status_im,
    input [6:0] io_cpu_ptw_status_zero,
    input  io_cpu_ptw_status_er,
    input  io_cpu_ptw_status_vm,
    input  io_cpu_ptw_status_s64,
    input  io_cpu_ptw_status_u64,
    input  io_cpu_ptw_status_ef,
    input  io_cpu_ptw_status_pei,
    input  io_cpu_ptw_status_ei,
    input  io_cpu_ptw_status_ps,
    input  io_cpu_ptw_status_s,
    input  io_cpu_ptw_invalidate,
    input  io_cpu_ptw_sret,
    output io_cpu_ordered,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[1:0] io_mem_acquire_bits_header_src,
    output[1:0] io_mem_acquire_bits_header_dst,
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[3:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [3:0] io_mem_grant_bits_payload_client_xact_id,
    input [3:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[3:0] io_mem_finish_bits_payload_master_xact_id,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [1:0] io_mem_probe_bits_header_src,
    input [1:0] io_mem_probe_bits_header_dst,
    input [25:0] io_mem_probe_bits_payload_addr,
    input [3:0] io_mem_probe_bits_payload_master_xact_id,
    input [1:0] io_mem_probe_bits_payload_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    output[1:0] io_mem_release_bits_header_src,
    output[1:0] io_mem_release_bits_header_dst,
    output[25:0] io_mem_release_bits_payload_addr,
    output[3:0] io_mem_release_bits_payload_client_xact_id,
    output[3:0] io_mem_release_bits_payload_master_xact_id,
    output[511:0] io_mem_release_bits_payload_data,
    output[2:0] io_mem_release_bits_payload_r_type
);

  wire wb_io_req_ready;
  wire[2:0] prober_io_wb_req_bits_r_type;
  wire[3:0] prober_io_wb_req_bits_master_xact_id;
  wire[3:0] prober_io_wb_req_bits_client_xact_id;
  wire prober_io_wb_req_bits_way_en;
  wire[5:0] prober_io_wb_req_bits_idx;
  wire[19:0] prober_io_wb_req_bits_tag;
  wire prober_io_wb_req_valid;
  wire[2:0] mshrs_io_wb_req_bits_r_type;
  wire[3:0] mshrs_io_wb_req_bits_master_xact_id;
  wire[3:0] mshrs_io_wb_req_bits_client_xact_id;
  wire mshrs_io_wb_req_bits_way_en;
  wire[5:0] mshrs_io_wb_req_bits_idx;
  wire[19:0] mshrs_io_wb_req_bits_tag;
  wire mshrs_io_wb_req_valid;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[3:0] FlowThroughSerializer_io_out_bits_payload_g_type;
  wire T4;
  wire writeArb_io_in_1_ready;
  wire T5;
  wire[2:0] wb_io_release_bits_r_type;
  wire[511:0] wb_io_release_bits_data;
  wire[3:0] wb_io_release_bits_master_xact_id;
  wire[3:0] wb_io_release_bits_client_xact_id;
  wire[25:0] wb_io_release_bits_addr;
  wire wb_io_release_valid;
  wire[2:0] prober_io_rep_bits_r_type;
  wire[511:0] prober_io_rep_bits_data;
  wire[3:0] prober_io_rep_bits_master_xact_id;
  wire[3:0] prober_io_rep_bits_client_xact_id;
  wire[25:0] prober_io_rep_bits_addr;
  wire prober_io_rep_valid;
  reg [63:0] s2_req_data;
  wire[63:0] T6;
  wire[63:0] T7;
  wire[63:0] T8;
  wire[63:0] mshrs_io_replay_bits_data;
  reg  s1_replay;
  wire T9;
  wire T10;
  wire readArb_io_in_1_ready;
  wire mshrs_io_replay_valid;
  wire T11;
  wire s1_write;
  wire T12;
  wire T13;
  reg [4:0] s1_req_cmd;
  wire[4:0] T14;
  wire[4:0] T15;
  wire[4:0] T16;
  wire[4:0] mshrs_io_replay_bits_cmd;
  reg [4:0] s2_req_cmd;
  wire[4:0] T17;
  reg  s1_clk_en;
  wire metaReadArb_io_out_valid;
  wire s2_recycle;
  wire T18;
  reg  s2_recycle_next;
  wire T19;
  wire T20;
  wire T21;
  wire s2_recycle_ecc;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  reg [43:0] s2_req_addr;
  wire[43:0] T28;
  wire[43:0] T29;
  wire[31:0] s1_addr;
  wire[12:0] T30;
  reg [43:0] s1_req_addr;
  wire[43:0] T31;
  wire[43:0] T32;
  wire[43:0] T33;
  wire[43:0] T34;
  wire[43:0] T35;
  wire[43:0] T36;
  wire[31:0] T37;
  wire[25:0] T38;
  wire[5:0] wb_io_meta_read_bits_idx;
  wire[19:0] wb_io_meta_read_bits_tag;
  wire wb_io_meta_read_valid;
  wire[43:0] T39;
  wire[31:0] T40;
  wire[25:0] T41;
  wire[5:0] prober_io_meta_read_bits_idx;
  wire[19:0] prober_io_meta_read_bits_tag;
  wire prober_io_meta_read_valid;
  wire[43:0] mshrs_io_replay_bits_addr;
  wire[18:0] dtlb_io_resp_ppn;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire s2_hit;
  wire T45;
  wire[1:0] T46;
  wire[1:0] T47;
  reg [1:0] s2_hit_state_state;
  wire[1:0] T48;
  wire[1:0] meta_io_resp_0_coh_state;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  reg  s2_tag_match_way;
  wire T78;
  wire s1_tag_match_way;
  wire T79;
  wire T80;
  wire T81;
  wire s1_tag_eq_way;
  wire T82;
  wire[19:0] T83;
  wire[19:0] meta_io_resp_0_tag;
  wire T84;
  wire s2_replay;
  wire T85;
  reg  R86;
  wire T87;
  reg  s2_valid;
  wire T88;
  wire s1_valid_masked;
  wire T89;
  reg  s1_valid;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  reg [63:0] s1_req_data;
  wire[63:0] T98;
  wire[63:0] T99;
  wire[63:0] T100;
  wire T101;
  reg  s1_recycled;
  wire T102;
  wire[63:0] T103;
  wire[127:0] s2_data_word;
  wire[127:0] s2_data_word_prebypass;
  wire[6:0] T104;
  wire[127:0] s2_data_uncorrected;
  wire[127:0] T105;
  wire[63:0] T106;
  wire[127:0] s2_data_muxed;
  wire[127:0] T107;
  wire[127:0] T108;
  reg [63:0] R109;
  wire[63:0] T110;
  wire[127:0] T111;
  wire[127:0] T112;
  wire[127:0] T113;
  wire[127:0] data_io_resp_0;
  wire T114;
  wire T115;
  reg [63:0] R116;
  wire[63:0] T117;
  wire[63:0] T118;
  wire[63:0] T119;
  wire[127:0] T120;
  reg [63:0] s2_store_bypass_data;
  wire[63:0] T121;
  wire[63:0] T122;
  wire[63:0] T123;
  reg [63:0] s4_req_data;
  wire[63:0] T124;
  reg [63:0] s3_req_data;
  wire[63:0] T125;
  wire[127:0] T126;
  wire[127:0] T127;
  wire[63:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire[127:0] T139;
  wire[127:0] T140;
  wire[63:0] amoalu_io_out;
  wire[127:0] s2_data_corrected;
  wire[127:0] T141;
  wire T142;
  reg  s3_valid;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire s2_sc_fail;
  wire T154;
  wire s2_lrsc_addr_match;
  wire T155;
  wire[37:0] T156;
  reg [37:0] lrsc_addr;
  wire[37:0] T157;
  wire[37:0] T158;
  wire T159;
  wire s2_lr;
  wire T160;
  wire T161;
  wire s2_valid_masked;
  wire T162;
  wire T163;
  wire s2_nack;
  wire s2_nack_miss;
  wire T164;
  wire mshrs_io_req_ready;
  wire T165;
  wire T166;
  wire s2_nack_victim;
  wire mshrs_io_secondary_miss;
  reg  s2_nack_hit;
  wire T167;
  wire s1_nack;
  wire T168;
  wire T169;
  wire prober_io_req_ready;
  wire T170;
  wire[5:0] prober_io_meta_write_bits_idx;
  wire[5:0] T171;
  wire T172;
  wire dtlb_io_resp_miss;
  wire T173;
  wire T174;
  reg [4:0] lrsc_count;
  wire[4:0] T175;
  wire[4:0] T176;
  wire[4:0] T177;
  wire[4:0] T178;
  wire[4:0] T179;
  wire[4:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire s2_sc;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  reg [4:0] s3_req_cmd;
  wire[4:0] T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[40:0] T197;
  reg [43:0] s3_req_addr;
  wire[43:0] T198;
  wire[40:0] T199;
  wire[28:0] T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire[40:0] T211;
  wire[40:0] T212;
  wire[28:0] T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  reg [4:0] s4_req_cmd;
  wire[4:0] T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire[40:0] T230;
  reg [43:0] s4_req_addr;
  wire[43:0] T231;
  wire[40:0] T232;
  wire[28:0] T233;
  reg  s4_valid;
  wire T234;
  wire T235;
  reg  s2_store_bypass;
  wire T236;
  wire T237;
  reg [2:0] s2_req_typ;
  wire[2:0] T238;
  reg [2:0] s1_req_typ;
  wire[2:0] T239;
  wire[2:0] T240;
  wire[2:0] T241;
  wire[2:0] mshrs_io_replay_bits_typ;
  wire[3:0] T242;
  wire[5:0] T243;
  wire data_io_write_ready;
  wire[127:0] T244;
  wire[1:0] T245;
  wire T246;
  wire T247;
  wire[11:0] T248;
  reg  s3_way;
  wire T249;
  wire[127:0] T250;
  wire[511:0] FlowThroughSerializer_io_out_bits_payload_data;
  wire[11:0] mshrs_io_mem_resp_addr;
  wire mshrs_io_mem_resp_way_en;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire FlowThroughSerializer_io_out_valid;
  wire T255;
  wire T256;
  wire[11:0] T257;
  wire[11:0] T258;
  wire[11:0] wb_io_data_req_bits_addr;
  wire wb_io_data_req_bits_way_en;
  wire wb_io_data_req_valid;
  wire[11:0] T259;
  wire[127:0] T260;
  wire[127:0] T261;
  wire[63:0] T262;
  wire[127:0] writeArb_io_out_bits_data;
  wire[63:0] T263;
  wire[1:0] writeArb_io_out_bits_wmask;
  wire[11:0] writeArb_io_out_bits_addr;
  wire writeArb_io_out_bits_way_en;
  wire writeArb_io_out_valid;
  wire[11:0] readArb_io_out_bits_addr;
  wire readArb_io_out_bits_way_en;
  wire readArb_io_out_valid;
  wire meta_io_write_ready;
  wire[1:0] mshrs_io_meta_write_bits_data_coh_state;
  wire[19:0] mshrs_io_meta_write_bits_data_tag;
  wire mshrs_io_meta_write_bits_way_en;
  wire[5:0] mshrs_io_meta_write_bits_idx;
  wire mshrs_io_meta_write_valid;
  wire[1:0] prober_io_meta_write_bits_data_coh_state;
  wire[19:0] prober_io_meta_write_bits_data_tag;
  wire prober_io_meta_write_bits_way_en;
  wire prober_io_meta_write_valid;
  wire meta_io_read_ready;
  wire[5:0] T264;
  wire[37:0] T265;
  wire[5:0] mshrs_io_meta_read_bits_idx;
  wire mshrs_io_meta_read_valid;
  wire[5:0] T266;
  wire[37:0] T267;
  wire[1:0] metaWriteArb_io_out_bits_data_coh_state;
  wire[19:0] metaWriteArb_io_out_bits_data_tag;
  wire metaWriteArb_io_out_bits_way_en;
  wire[5:0] metaWriteArb_io_out_bits_idx;
  wire metaWriteArb_io_out_valid;
  wire[5:0] metaReadArb_io_out_bits_idx;
  reg  s1_req_phys;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire mshrs_io_replay_bits_phys;
  reg  s2_req_phys;
  wire T273;
  wire[30:0] T274;
  wire T275;
  wire T276;
  wire T277;
  wire s1_readwrite;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire s1_read;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire wbArb_io_in_1_ready;
  wire[3:0] FlowThroughSerializer_io_out_bits_payload_master_xact_id;
  wire[3:0] FlowThroughSerializer_io_out_bits_payload_client_xact_id;
  wire[1:0] FlowThroughSerializer_io_out_bits_header_dst;
  wire[1:0] FlowThroughSerializer_io_out_bits_header_src;
  wire T288;
  wire metaWriteArb_io_in_0_ready;
  wire metaReadArb_io_in_1_ready;
  wire T289;
  wire T290;
  wire[1:0] T291;
  wire[1:0] s2_replaced_way_en;
  reg  R292;
  wire T293;
  wire[1:0] T294;
  wire[1:0] T295;
  wire[21:0] T296;
  wire[21:0] T297;
  reg [1:0] s2_repl_meta_coh_state;
  wire[1:0] T298;
  reg [19:0] s2_repl_meta_tag;
  wire[19:0] T299;
  wire[21:0] T300;
  wire[1:0] T301;
  wire[19:0] T302;
  wire[19:0] T303;
  reg [7:0] s2_req_tag;
  wire[7:0] T304;
  reg [7:0] s1_req_tag;
  wire[7:0] T305;
  wire[7:0] T306;
  wire[7:0] T307;
  wire[7:0] mshrs_io_replay_bits_tag;
  reg  s2_req_kill;
  wire T308;
  reg  s1_req_kill;
  wire T309;
  wire T310;
  wire T311;
  wire mshrs_io_replay_bits_kill;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire mshrs_io_probe_rdy;
  wire wbArb_io_in_0_ready;
  wire metaWriteArb_io_in_1_ready;
  wire metaReadArb_io_in_2_ready;
  wire releaseArb_io_in_1_ready;
  wire[1:0] probe_bits_p_type;
  wire[3:0] probe_bits_master_xact_id;
  wire[25:0] probe_bits_addr;
  wire T335;
  wire T336;
  wire probe_valid;
  wire releaseArb_io_in_0_ready;
  wire readArb_io_in_2_ready;
  wire metaReadArb_io_in_3_ready;
  wire[2:0] wbArb_io_out_bits_r_type;
  wire[3:0] wbArb_io_out_bits_master_xact_id;
  wire[3:0] wbArb_io_out_bits_client_xact_id;
  wire wbArb_io_out_bits_way_en;
  wire[5:0] wbArb_io_out_bits_idx;
  wire[19:0] wbArb_io_out_bits_tag;
  wire wbArb_io_out_valid;
  wire[2:0] T337;
  wire[2:0] releaseArb_io_out_bits_r_type;
  wire[511:0] T338;
  wire[511:0] releaseArb_io_out_bits_data;
  wire[3:0] T339;
  wire[3:0] releaseArb_io_out_bits_master_xact_id;
  wire[3:0] T340;
  wire[3:0] releaseArb_io_out_bits_client_xact_id;
  wire[25:0] T341;
  wire[25:0] releaseArb_io_out_bits_addr;
  wire[1:0] T342;
  wire[1:0] T343;
  wire T344;
  wire releaseArb_io_out_valid;
  wire probe_ready;
  wire T345;
  wire T346;
  wire[3:0] mshrs_io_mem_finish_bits_payload_master_xact_id;
  wire[1:0] mshrs_io_mem_finish_bits_header_dst;
  wire[1:0] mshrs_io_mem_finish_bits_header_src;
  wire mshrs_io_mem_finish_valid;
  wire FlowThroughSerializer_io_in_ready;
  wire[3:0] T347;
  wire[3:0] mshrs_io_mem_req_bits_atomic_opcode;
  wire[2:0] T348;
  wire[2:0] mshrs_io_mem_req_bits_subword_addr;
  wire[5:0] T349;
  wire[5:0] mshrs_io_mem_req_bits_write_mask;
  wire[2:0] T350;
  wire[2:0] mshrs_io_mem_req_bits_a_type;
  wire[511:0] T351;
  wire[511:0] mshrs_io_mem_req_bits_data;
  wire[3:0] T352;
  wire[3:0] mshrs_io_mem_req_bits_client_xact_id;
  wire[25:0] T353;
  wire[25:0] mshrs_io_mem_req_bits_addr;
  wire[1:0] T354;
  wire[1:0] T355;
  wire T356;
  wire mshrs_io_mem_req_valid;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire mshrs_io_fence_rdy;
  wire[29:0] dtlb_io_ptw_req_bits;
  wire dtlb_io_ptw_req_valid;
  wire T361;
  wire dtlb_io_resp_xcpt_st;
  wire T362;
  wire dtlb_io_resp_xcpt_ld;
  wire T363;
  wire misaligned;
  wire T364;
  wire T365;
  wire[2:0] T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire[1:0] T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire s1_sc;
  wire[3:0] T384;
  wire[63:0] T385;
  wire[63:0] T386;
  wire[63:0] T387;
  wire[7:0] T388;
  wire[7:0] T389;
  wire[7:0] T390;
  wire[63:0] T391;
  wire[15:0] T392;
  wire[15:0] T393;
  wire[63:0] T394;
  wire[31:0] T395;
  wire[31:0] T396;
  wire[31:0] T397;
  wire T398;
  wire[31:0] T399;
  wire[31:0] T400;
  wire[31:0] T401;
  wire[31:0] T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire[15:0] T415;
  wire T416;
  wire[47:0] T417;
  wire[47:0] T418;
  wire[47:0] T419;
  wire[47:0] T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire[7:0] T426;
  wire T427;
  wire[55:0] T428;
  wire[55:0] T429;
  wire[55:0] T430;
  wire[55:0] T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire dtlb_io_req_ready;
  wire T458;
  wire metaReadArb_io_in_4_ready;
  wire T459;
  wire readArb_io_in_3_ready;
  reg  block_miss;
  wire T460;
  wire T461;
  wire T462;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    s2_req_data = {2{$random}};
    s1_replay = {1{$random}};
    s1_req_cmd = {1{$random}};
    s2_req_cmd = {1{$random}};
    s1_clk_en = {1{$random}};
    s2_recycle_next = {1{$random}};
    s2_req_addr = {2{$random}};
    s1_req_addr = {2{$random}};
    s2_hit_state_state = {1{$random}};
    s2_tag_match_way = {1{$random}};
    R86 = {1{$random}};
    s2_valid = {1{$random}};
    s1_valid = {1{$random}};
    s1_req_data = {2{$random}};
    s1_recycled = {1{$random}};
    R109 = {2{$random}};
    R116 = {2{$random}};
    s2_store_bypass_data = {2{$random}};
    s4_req_data = {2{$random}};
    s3_req_data = {2{$random}};
    s3_valid = {1{$random}};
    lrsc_addr = {2{$random}};
    s2_nack_hit = {1{$random}};
    lrsc_count = {1{$random}};
    s3_req_cmd = {1{$random}};
    s3_req_addr = {2{$random}};
    s4_req_cmd = {1{$random}};
    s4_req_addr = {2{$random}};
    s4_valid = {1{$random}};
    s2_store_bypass = {1{$random}};
    s2_req_typ = {1{$random}};
    s1_req_typ = {1{$random}};
    s3_way = {1{$random}};
    s1_req_phys = {1{$random}};
    s2_req_phys = {1{$random}};
    R292 = {1{$random}};
    s2_repl_meta_coh_state = {1{$random}};
    s2_repl_meta_tag = {1{$random}};
    s2_req_tag = {1{$random}};
    s1_req_tag = {1{$random}};
    s2_req_kill = {1{$random}};
    s1_req_kill = {1{$random}};
    block_miss = {1{$random}};
  end
`endif

  assign T0 = writeArb_io_in_1_ready | T1;
  assign T1 = T2 ^ 1'h1;
  assign T2 = T4 | T3;
  assign T3 = FlowThroughSerializer_io_out_bits_payload_g_type == 4'h2;
  assign T4 = FlowThroughSerializer_io_out_bits_payload_g_type == 4'h1;
  assign T5 = io_mem_release_ready;
  assign T6 = T101 ? s1_req_data : T7;
  assign T7 = T11 ? T8 : s2_req_data;
  assign T8 = s1_replay ? mshrs_io_replay_bits_data : io_cpu_req_bits_data;
  assign T9 = reset ? 1'h0 : T10;
  assign T10 = mshrs_io_replay_valid & readArb_io_in_1_ready;
  assign T11 = s1_clk_en & s1_write;
  assign s1_write = T95 | T12;
  assign T12 = T94 | T13;
  assign T13 = s1_req_cmd == 5'h4;
  assign T14 = s2_recycle ? s2_req_cmd : T15;
  assign T15 = mshrs_io_replay_valid ? mshrs_io_replay_bits_cmd : T16;
  assign T16 = io_cpu_req_valid ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign T17 = s1_clk_en ? s1_req_cmd : s2_req_cmd;
  assign s2_recycle = T18;
  assign T18 = s2_recycle_ecc | s2_recycle_next;
  assign T19 = reset ? 1'h0 : T20;
  assign T20 = T93 ? T21 : s2_recycle_next;
  assign T21 = T92 & s2_recycle_ecc;
  assign s2_recycle_ecc = T44 & T22;
  assign T22 = T42 & T23;
  assign T23 = T24 - 1'h1;
  assign T24 = 1'h1 << T25;
  assign T25 = T26 + 1'h1;
  assign T26 = T27 - T27;
  assign T27 = s2_req_addr[2'h3:2'h3];
  assign T28 = s1_clk_en ? T29 : s2_req_addr;
  assign T29 = {12'h0, s1_addr};
  assign s1_addr = {dtlb_io_resp_ppn, T30};
  assign T30 = s1_req_addr[4'hc:1'h0];
  assign T31 = s2_recycle ? s2_req_addr : T32;
  assign T32 = mshrs_io_replay_valid ? mshrs_io_replay_bits_addr : T33;
  assign T33 = prober_io_meta_read_valid ? T39 : T34;
  assign T34 = wb_io_meta_read_valid ? T36 : T35;
  assign T35 = io_cpu_req_valid ? io_cpu_req_bits_addr : s1_req_addr;
  assign T36 = {12'h0, T37};
  assign T37 = T38 << 3'h6;
  assign T38 = {wb_io_meta_read_bits_tag, wb_io_meta_read_bits_idx};
  assign T39 = {12'h0, T40};
  assign T40 = T41 << 3'h6;
  assign T41 = {prober_io_meta_read_bits_tag, prober_io_meta_read_bits_idx};
  assign T42 = T43 >> T27;
  assign T43 = 2'h0;
  assign T44 = T84 & s2_hit;
  assign s2_hit = T56 & T45;
  assign T45 = s2_hit_state_state == T46;
  assign T46 = T47;
  assign T47 = T49 ? 2'h3 : s2_hit_state_state;
  assign T48 = s1_clk_en ? meta_io_resp_0_coh_state : s2_hit_state_state;
  assign T49 = T53 | T50;
  assign T50 = T52 | T51;
  assign T51 = s2_req_cmd == 5'h4;
  assign T52 = s2_req_cmd[2'h3:2'h3];
  assign T53 = T55 | T54;
  assign T54 = s2_req_cmd == 5'h7;
  assign T55 = s2_req_cmd == 5'h1;
  assign T56 = T77 & T57;
  assign T57 = T66 ? T63 : T58;
  assign T58 = T60 | T59;
  assign T59 = s2_hit_state_state == 2'h3;
  assign T60 = T62 | T61;
  assign T61 = s2_hit_state_state == 2'h2;
  assign T62 = s2_hit_state_state == 2'h1;
  assign T63 = T65 | T64;
  assign T64 = s2_hit_state_state == 2'h3;
  assign T65 = s2_hit_state_state == 2'h2;
  assign T66 = T68 | T67;
  assign T67 = s2_req_cmd == 5'h6;
  assign T68 = T70 | T69;
  assign T69 = s2_req_cmd == 5'h3;
  assign T70 = T74 | T71;
  assign T71 = T73 | T72;
  assign T72 = s2_req_cmd == 5'h4;
  assign T73 = s2_req_cmd[2'h3:2'h3];
  assign T74 = T76 | T75;
  assign T75 = s2_req_cmd == 5'h7;
  assign T76 = s2_req_cmd == 5'h1;
  assign T77 = s2_tag_match_way != 1'h0;
  assign T78 = s1_clk_en ? s1_tag_match_way : s2_tag_match_way;
  assign s1_tag_match_way = T79;
  assign T79 = T81 & T80;
  assign T80 = meta_io_resp_0_coh_state != 2'h0;
  assign T81 = s1_tag_eq_way;
  assign s1_tag_eq_way = T82;
  assign T82 = meta_io_resp_0_tag == T83;
  assign T83 = s1_addr >> 4'hc;
  assign T84 = s2_valid | s2_replay;
  assign s2_replay = R86 & T85;
  assign T85 = s2_req_cmd != 5'h5;
  assign T87 = reset ? 1'h0 : s1_replay;
  assign T88 = reset ? 1'h0 : s1_valid_masked;
  assign s1_valid_masked = s1_valid & T89;
  assign T89 = io_cpu_req_bits_kill ^ 1'h1;
  assign T90 = reset ? 1'h0 : T91;
  assign T91 = io_cpu_req_ready & io_cpu_req_valid;
  assign T92 = s1_valid | s1_replay;
  assign T93 = s1_valid | s1_replay;
  assign T94 = s1_req_cmd[2'h3:2'h3];
  assign T95 = T97 | T96;
  assign T96 = s1_req_cmd == 5'h7;
  assign T97 = s1_req_cmd == 5'h1;
  assign T98 = s2_recycle ? s2_req_data : T99;
  assign T99 = mshrs_io_replay_valid ? mshrs_io_replay_bits_data : T100;
  assign T100 = io_cpu_req_valid ? io_cpu_req_bits_data : s1_req_data;
  assign T101 = s1_clk_en & s1_recycled;
  assign T102 = s1_clk_en ? s2_recycle : s1_recycled;
  assign T103 = s2_data_word[6'h3f:1'h0];
  assign s2_data_word = s2_store_bypass ? T120 : s2_data_word_prebypass;
  assign s2_data_word_prebypass = s2_data_uncorrected >> T104;
  assign T104 = {T27, 6'h0};
  assign s2_data_uncorrected = T105;
  assign T105 = {T119, T106};
  assign T106 = s2_data_muxed[6'h3f:1'h0];
  assign s2_data_muxed = T107;
  assign T107 = T108;
  assign T108 = {R116, R109};
  assign T110 = T111[6'h3f:1'h0];
  assign T111 = T114 ? T113 : T112;
  assign T112 = {64'h0, R109};
  assign T113 = data_io_resp_0 >> 1'h0;
  assign T114 = s1_clk_en & T115;
  assign T115 = s1_tag_eq_way;
  assign T117 = T114 ? T118 : R116;
  assign T118 = data_io_resp_0 >> 7'h40;
  assign T119 = s2_data_muxed[7'h7f:7'h40];
  assign T120 = {64'h0, s2_store_bypass_data};
  assign T121 = T217 ? T122 : s2_store_bypass_data;
  assign T122 = T201 ? amoalu_io_out : T123;
  assign T123 = T186 ? s3_req_data : s4_req_data;
  assign T124 = T142 ? s3_req_data : s4_req_data;
  assign T125 = T126[6'h3f:1'h0];
  assign T126 = T129 ? T139 : T127;
  assign T127 = {64'h0, T128};
  assign T128 = T129 ? s2_req_data : s3_req_data;
  assign T129 = T138 & T130;
  assign T130 = T131 | T22;
  assign T131 = T135 | T132;
  assign T132 = T134 | T133;
  assign T133 = s2_req_cmd == 5'h4;
  assign T134 = s2_req_cmd[2'h3:2'h3];
  assign T135 = T137 | T136;
  assign T136 = s2_req_cmd == 5'h7;
  assign T137 = s2_req_cmd == 5'h1;
  assign T138 = s2_valid | s2_replay;
  assign T139 = T22 ? s2_data_corrected : T140;
  assign T140 = {64'h0, amoalu_io_out};
  assign s2_data_corrected = T141;
  assign T141 = {T119, T106};
  assign T142 = s3_valid & metaReadArb_io_out_valid;
  assign T143 = reset ? 1'h0 : T144;
  assign T144 = T152 & T145;
  assign T145 = T149 | T146;
  assign T146 = T148 | T147;
  assign T147 = s2_req_cmd == 5'h4;
  assign T148 = s2_req_cmd[2'h3:2'h3];
  assign T149 = T151 | T150;
  assign T150 = s2_req_cmd == 5'h7;
  assign T151 = s2_req_cmd == 5'h1;
  assign T152 = T184 & T153;
  assign T153 = s2_sc_fail ^ 1'h1;
  assign s2_sc_fail = s2_sc & T154;
  assign T154 = s2_lrsc_addr_match ^ 1'h1;
  assign s2_lrsc_addr_match = T174 & T155;
  assign T155 = lrsc_addr == T156;
  assign T156 = s2_req_addr >> 3'h6;
  assign T157 = T159 ? T158 : lrsc_addr;
  assign T158 = s2_req_addr >> 3'h6;
  assign T159 = T160 & s2_lr;
  assign s2_lr = s2_req_cmd == 5'h6;
  assign T160 = T161 | s2_replay;
  assign T161 = s2_valid_masked & s2_hit;
  assign s2_valid_masked = T162;
  assign T162 = s2_valid & T163;
  assign T163 = s2_nack ^ 1'h1;
  assign s2_nack = T166 | s2_nack_miss;
  assign s2_nack_miss = T165 & T164;
  assign T164 = mshrs_io_req_ready ^ 1'h1;
  assign T165 = s2_hit ^ 1'h1;
  assign T166 = s2_nack_hit | s2_nack_victim;
  assign s2_nack_victim = s2_hit & mshrs_io_secondary_miss;
  assign T167 = T173 ? s1_nack : s2_nack_hit;
  assign s1_nack = T172 | T168;
  assign T168 = T170 & T169;
  assign T169 = prober_io_req_ready ^ 1'h1;
  assign T170 = T171 == prober_io_meta_write_bits_idx;
  assign T171 = s1_req_addr[4'hb:3'h6];
  assign T172 = T275 & dtlb_io_resp_miss;
  assign T173 = s1_valid | s1_replay;
  assign T174 = lrsc_count != 5'h0;
  assign T175 = reset ? 5'h0 : T176;
  assign T176 = io_cpu_ptw_sret ? 5'h0 : T177;
  assign T177 = T183 ? 5'h0 : T178;
  assign T178 = T181 ? 5'h1f : T179;
  assign T179 = T174 ? T180 : lrsc_count;
  assign T180 = lrsc_count - 5'h1;
  assign T181 = T159 & T182;
  assign T182 = T174 ^ 1'h1;
  assign T183 = T160 & s2_sc;
  assign s2_sc = s2_req_cmd == 5'h7;
  assign T184 = T185 | s2_replay;
  assign T185 = s2_valid_masked & s2_hit;
  assign T186 = T195 & T187;
  assign T187 = T192 | T188;
  assign T188 = T191 | T189;
  assign T189 = s3_req_cmd == 5'h4;
  assign T190 = T129 ? s2_req_cmd : s3_req_cmd;
  assign T191 = s3_req_cmd[2'h3:2'h3];
  assign T192 = T194 | T193;
  assign T193 = s3_req_cmd == 5'h7;
  assign T194 = s3_req_cmd == 5'h1;
  assign T195 = s3_valid & T196;
  assign T196 = T199 == T197;
  assign T197 = s3_req_addr >> 2'h3;
  assign T198 = T129 ? s2_req_addr : s3_req_addr;
  assign T199 = {12'h0, T200};
  assign T200 = s1_addr >> 2'h3;
  assign T201 = T209 & T202;
  assign T202 = T206 | T203;
  assign T203 = T205 | T204;
  assign T204 = s2_req_cmd == 5'h4;
  assign T205 = s2_req_cmd[2'h3:2'h3];
  assign T206 = T208 | T207;
  assign T207 = s2_req_cmd == 5'h7;
  assign T208 = s2_req_cmd == 5'h1;
  assign T209 = T214 & T210;
  assign T210 = T212 == T211;
  assign T211 = s2_req_addr >> 2'h3;
  assign T212 = {12'h0, T213};
  assign T213 = s1_addr >> 2'h3;
  assign T214 = T216 & T215;
  assign T215 = s2_sc_fail ^ 1'h1;
  assign T216 = s2_valid_masked | s2_replay;
  assign T217 = s1_clk_en & T218;
  assign T218 = T235 | T219;
  assign T219 = T228 & T220;
  assign T220 = T225 | T221;
  assign T221 = T224 | T222;
  assign T222 = s4_req_cmd == 5'h4;
  assign T223 = T142 ? s3_req_cmd : s4_req_cmd;
  assign T224 = s4_req_cmd[2'h3:2'h3];
  assign T225 = T227 | T226;
  assign T226 = s4_req_cmd == 5'h7;
  assign T227 = s4_req_cmd == 5'h1;
  assign T228 = s4_valid & T229;
  assign T229 = T232 == T230;
  assign T230 = s4_req_addr >> 2'h3;
  assign T231 = T142 ? s3_req_addr : s4_req_addr;
  assign T232 = {12'h0, T233};
  assign T233 = s1_addr >> 2'h3;
  assign T234 = reset ? 1'h0 : s3_valid;
  assign T235 = T201 | T186;
  assign T236 = T217 ? 1'h1 : T237;
  assign T237 = s1_clk_en ? 1'h0 : s2_store_bypass;
  assign T238 = s1_clk_en ? s1_req_typ : s2_req_typ;
  assign T239 = s2_recycle ? s2_req_typ : T240;
  assign T240 = mshrs_io_replay_valid ? mshrs_io_replay_bits_typ : T241;
  assign T241 = io_cpu_req_valid ? io_cpu_req_bits_typ : s1_req_typ;
  assign T242 = s2_req_cmd[2'h3:1'h0];
  assign T243 = s2_req_addr[3'h5:1'h0];
  assign T244 = {s3_req_data, s3_req_data};
  assign T245 = 1'h1 << T246;
  assign T246 = T247;
  assign T247 = s3_req_addr[2'h3:2'h3];
  assign T248 = s3_req_addr[4'hb:1'h0];
  assign T249 = T129 ? s2_tag_match_way : s3_way;
  assign T250 = FlowThroughSerializer_io_out_bits_payload_data[7'h7f:1'h0];
  assign T251 = FlowThroughSerializer_io_out_valid & T252;
  assign T252 = T254 | T253;
  assign T253 = FlowThroughSerializer_io_out_bits_payload_g_type == 4'h2;
  assign T254 = FlowThroughSerializer_io_out_bits_payload_g_type == 4'h1;
  assign T255 = T256 | T0;
  assign T256 = FlowThroughSerializer_io_out_valid ^ 1'h1;
  assign T257 = s2_req_addr[4'hb:1'h0];
  assign T258 = mshrs_io_replay_bits_addr[4'hb:1'h0];
  assign T259 = io_cpu_req_bits_addr[4'hb:1'h0];
  assign T260 = T261;
  assign T261 = {T263, T262};
  assign T262 = writeArb_io_out_bits_data[6'h3f:1'h0];
  assign T263 = writeArb_io_out_bits_data[7'h7f:7'h40];
  assign T264 = T265[3'h5:1'h0];
  assign T265 = s2_req_addr >> 3'h6;
  assign T266 = T267[3'h5:1'h0];
  assign T267 = io_cpu_req_bits_addr >> 3'h6;
  assign T268 = s2_recycle ? s2_req_phys : T269;
  assign T269 = mshrs_io_replay_valid ? mshrs_io_replay_bits_phys : T270;
  assign T270 = prober_io_meta_read_valid ? 1'h1 : T271;
  assign T271 = wb_io_meta_read_valid ? 1'h1 : T272;
  assign T272 = io_cpu_req_valid ? io_cpu_req_bits_phys : s1_req_phys;
  assign T273 = s1_clk_en ? s1_req_phys : s2_req_phys;
  assign T274 = s1_req_addr >> 4'hd;
  assign T275 = T277 & T276;
  assign T276 = s1_req_phys ^ 1'h1;
  assign T277 = s1_valid_masked & s1_readwrite;
  assign s1_readwrite = T281 | T278;
  assign T278 = T280 | T279;
  assign T279 = s1_req_cmd == 5'h3;
  assign T280 = s1_req_cmd == 5'h2;
  assign T281 = s1_read | s1_write;
  assign s1_read = T285 | T282;
  assign T282 = T284 | T283;
  assign T283 = s1_req_cmd == 5'h4;
  assign T284 = s1_req_cmd[2'h3:2'h3];
  assign T285 = T287 | T286;
  assign T286 = s1_req_cmd == 5'h6;
  assign T287 = s1_req_cmd == 5'h0;
  assign T288 = T0 & FlowThroughSerializer_io_out_valid;
  assign T289 = io_mem_acquire_ready;
  assign T290 = T291[1'h0:1'h0];
  assign T291 = T77 ? T294 : s2_replaced_way_en;
  assign s2_replaced_way_en = 1'h1 << R292;
  assign T293 = s1_clk_en ? 1'h0 : R292;
  assign T294 = {1'h0, s2_tag_match_way};
  assign T295 = T296[1'h1:1'h0];
  assign T296 = T77 ? T300 : T297;
  assign T297 = {s2_repl_meta_tag, s2_repl_meta_coh_state};
  assign T298 = s1_clk_en ? meta_io_resp_0_coh_state : s2_repl_meta_coh_state;
  assign T299 = s1_clk_en ? meta_io_resp_0_tag : s2_repl_meta_tag;
  assign T300 = {T302, T301};
  assign T301 = s2_hit_state_state;
  assign T302 = s2_repl_meta_tag;
  assign T303 = T296[5'h15:2'h2];
  assign T304 = s1_clk_en ? s1_req_tag : s2_req_tag;
  assign T305 = s2_recycle ? s2_req_tag : T306;
  assign T306 = mshrs_io_replay_valid ? mshrs_io_replay_bits_tag : T307;
  assign T307 = io_cpu_req_valid ? io_cpu_req_bits_tag : s1_req_tag;
  assign T308 = s1_clk_en ? s1_req_kill : s2_req_kill;
  assign T309 = s2_recycle ? s2_req_kill : T310;
  assign T310 = mshrs_io_replay_valid ? mshrs_io_replay_bits_kill : T311;
  assign T311 = io_cpu_req_valid ? io_cpu_req_bits_kill : s1_req_kill;
  assign T312 = s2_nack_hit ? 1'h0 : T313;
  assign T313 = T333 & T314;
  assign T314 = T322 | T315;
  assign T315 = T319 | T316;
  assign T316 = T318 | T317;
  assign T317 = s2_req_cmd == 5'h4;
  assign T318 = s2_req_cmd[2'h3:2'h3];
  assign T319 = T321 | T320;
  assign T320 = s2_req_cmd == 5'h7;
  assign T321 = s2_req_cmd == 5'h1;
  assign T322 = T330 | T323;
  assign T323 = T327 | T324;
  assign T324 = T326 | T325;
  assign T325 = s2_req_cmd == 5'h4;
  assign T326 = s2_req_cmd[2'h3:2'h3];
  assign T327 = T329 | T328;
  assign T328 = s2_req_cmd == 5'h6;
  assign T329 = s2_req_cmd == 5'h0;
  assign T330 = T332 | T331;
  assign T331 = s2_req_cmd == 5'h3;
  assign T332 = s2_req_cmd == 5'h2;
  assign T333 = s2_valid_masked & T334;
  assign T334 = s2_hit ^ 1'h1;
  assign probe_bits_p_type = io_mem_probe_bits_payload_p_type;
  assign probe_bits_master_xact_id = io_mem_probe_bits_payload_master_xact_id;
  assign probe_bits_addr = io_mem_probe_bits_payload_addr;
  assign T335 = probe_valid & T336;
  assign T336 = T174 ^ 1'h1;
  assign probe_valid = io_mem_probe_valid;
  assign io_mem_release_bits_payload_r_type = T337;
  assign T337 = releaseArb_io_out_bits_r_type;
  assign io_mem_release_bits_payload_data = T338;
  assign T338 = releaseArb_io_out_bits_data;
  assign io_mem_release_bits_payload_master_xact_id = T339;
  assign T339 = releaseArb_io_out_bits_master_xact_id;
  assign io_mem_release_bits_payload_client_xact_id = T340;
  assign T340 = releaseArb_io_out_bits_client_xact_id;
  assign io_mem_release_bits_payload_addr = T341;
  assign T341 = releaseArb_io_out_bits_addr;
  assign io_mem_release_bits_header_dst = T342;
  assign T342 = 2'h0;
  assign io_mem_release_bits_header_src = T343;
  assign T343 = 2'h0;
  assign io_mem_release_valid = T344;
  assign T344 = releaseArb_io_out_valid;
  assign io_mem_probe_ready = probe_ready;
  assign probe_ready = T345;
  assign T345 = prober_io_req_ready & T346;
  assign T346 = T174 ^ 1'h1;
  assign io_mem_finish_bits_payload_master_xact_id = mshrs_io_mem_finish_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = mshrs_io_mem_finish_bits_header_dst;
  assign io_mem_finish_bits_header_src = mshrs_io_mem_finish_bits_header_src;
  assign io_mem_finish_valid = mshrs_io_mem_finish_valid;
  assign io_mem_grant_ready = FlowThroughSerializer_io_in_ready;
  assign io_mem_acquire_bits_payload_atomic_opcode = T347;
  assign T347 = mshrs_io_mem_req_bits_atomic_opcode;
  assign io_mem_acquire_bits_payload_subword_addr = T348;
  assign T348 = mshrs_io_mem_req_bits_subword_addr;
  assign io_mem_acquire_bits_payload_write_mask = T349;
  assign T349 = mshrs_io_mem_req_bits_write_mask;
  assign io_mem_acquire_bits_payload_a_type = T350;
  assign T350 = mshrs_io_mem_req_bits_a_type;
  assign io_mem_acquire_bits_payload_data = T351;
  assign T351 = mshrs_io_mem_req_bits_data;
  assign io_mem_acquire_bits_payload_client_xact_id = T352;
  assign T352 = mshrs_io_mem_req_bits_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = T353;
  assign T353 = mshrs_io_mem_req_bits_addr;
  assign io_mem_acquire_bits_header_dst = T354;
  assign T354 = 2'h0;
  assign io_mem_acquire_bits_header_src = T355;
  assign T355 = 2'h0;
  assign io_mem_acquire_valid = T356;
  assign T356 = mshrs_io_mem_req_valid;
  assign io_cpu_ordered = T357;
  assign T357 = T359 & T358;
  assign T358 = s2_valid ^ 1'h1;
  assign T359 = mshrs_io_fence_rdy & T360;
  assign T360 = s1_valid ^ 1'h1;
  assign io_cpu_ptw_req_bits = dtlb_io_ptw_req_bits;
  assign io_cpu_ptw_req_valid = dtlb_io_ptw_req_valid;
  assign io_cpu_xcpt_pf_st = T361;
  assign T361 = s1_write & dtlb_io_resp_xcpt_st;
  assign io_cpu_xcpt_pf_ld = T362;
  assign T362 = s1_read & dtlb_io_resp_xcpt_ld;
  assign io_cpu_xcpt_ma_st = T363;
  assign T363 = s1_write & misaligned;
  assign misaligned = T368 | T364;
  assign T364 = T367 & T365;
  assign T365 = T366 != 3'h0;
  assign T366 = s1_req_addr[2'h2:1'h0];
  assign T367 = s1_req_typ == 3'h3;
  assign T368 = T375 | T369;
  assign T369 = T372 & T370;
  assign T370 = T371 != 2'h0;
  assign T371 = s1_req_addr[1'h1:1'h0];
  assign T372 = T374 | T373;
  assign T373 = s1_req_typ == 3'h6;
  assign T374 = s1_req_typ == 3'h2;
  assign T375 = T378 & T376;
  assign T376 = T377 != 1'h0;
  assign T377 = s1_req_addr[1'h0:1'h0];
  assign T378 = T380 | T379;
  assign T379 = s1_req_typ == 3'h5;
  assign T380 = s1_req_typ == 3'h1;
  assign io_cpu_xcpt_ma_ld = T381;
  assign T381 = s1_read & misaligned;
  assign io_cpu_replay_next_bits = s1_req_tag;
  assign io_cpu_replay_next_valid = T382;
  assign T382 = s1_replay & T383;
  assign T383 = s1_read | s1_sc;
  assign s1_sc = s1_req_cmd == 5'h7;
  assign io_cpu_resp_bits_store_data = s2_req_data;
  assign io_cpu_resp_bits_addr = s2_req_addr;
  assign io_cpu_resp_bits_cmd = T384;
  assign T384 = s2_req_cmd[2'h3:1'h0];
  assign io_cpu_resp_bits_tag = s2_req_tag;
  assign io_cpu_resp_bits_data_subword = T385;
  assign T385 = T387 | T386;
  assign T386 = {63'h0, s2_sc_fail};
  assign T387 = {T428, T388};
  assign T388 = s2_sc ? 8'h0 : T389;
  assign T389 = T427 ? T426 : T390;
  assign T390 = T391[3'h7:1'h0];
  assign T391 = {T417, T392};
  assign T392 = T416 ? T415 : T393;
  assign T393 = T394[4'hf:1'h0];
  assign T394 = {T399, T395};
  assign T395 = T398 ? T397 : T396;
  assign T396 = s2_data_word[5'h1f:1'h0];
  assign T397 = s2_data_word[6'h3f:6'h20];
  assign T398 = s2_req_addr[2'h2:2'h2];
  assign T399 = T412 ? T401 : T400;
  assign T400 = s2_data_word[6'h3f:6'h20];
  assign T401 = 32'h0 - T402;
  assign T402 = {31'h0, T403};
  assign T403 = T405 & T404;
  assign T404 = T395[5'h1f:5'h1f];
  assign T405 = T407 | T406;
  assign T406 = s2_req_typ == 3'h3;
  assign T407 = T409 | T408;
  assign T408 = s2_req_typ == 3'h2;
  assign T409 = T411 | T410;
  assign T410 = s2_req_typ == 3'h1;
  assign T411 = s2_req_typ == 3'h0;
  assign T412 = T414 | T413;
  assign T413 = s2_req_typ == 3'h6;
  assign T414 = s2_req_typ == 3'h2;
  assign T415 = T394[5'h1f:5'h10];
  assign T416 = s2_req_addr[1'h1:1'h1];
  assign T417 = T423 ? T419 : T418;
  assign T418 = T394[6'h3f:5'h10];
  assign T419 = 48'h0 - T420;
  assign T420 = {47'h0, T421};
  assign T421 = T405 & T422;
  assign T422 = T392[4'hf:4'hf];
  assign T423 = T425 | T424;
  assign T424 = s2_req_typ == 3'h5;
  assign T425 = s2_req_typ == 3'h1;
  assign T426 = T391[4'hf:4'h8];
  assign T427 = s2_req_addr[1'h0:1'h0];
  assign T428 = T434 ? T430 : T429;
  assign T429 = T391[6'h3f:4'h8];
  assign T430 = 56'h0 - T431;
  assign T431 = {55'h0, T432};
  assign T432 = T405 & T433;
  assign T433 = T388[3'h7:3'h7];
  assign T434 = s2_sc | T435;
  assign T435 = T437 | T436;
  assign T436 = s2_req_typ == 3'h4;
  assign T437 = s2_req_typ == 3'h0;
  assign io_cpu_resp_bits_data = T394;
  assign io_cpu_resp_bits_has_data = T438;
  assign T438 = T439 | s2_sc;
  assign T439 = T443 | T440;
  assign T440 = T442 | T441;
  assign T441 = s2_req_cmd == 5'h4;
  assign T442 = s2_req_cmd[2'h3:2'h3];
  assign T443 = T445 | T444;
  assign T444 = s2_req_cmd == 5'h6;
  assign T445 = s2_req_cmd == 5'h0;
  assign io_cpu_resp_bits_typ = s2_req_typ;
  assign io_cpu_resp_bits_replay = s2_replay;
  assign io_cpu_resp_bits_nack = T446;
  assign T446 = s2_valid & s2_nack;
  assign io_cpu_resp_valid = T447;
  assign T447 = T449 & T448;
  assign T448 = T22 ^ 1'h1;
  assign T449 = s2_replay | T450;
  assign T450 = s2_valid_masked & s2_hit;
  assign io_cpu_req_ready = T451;
  assign T451 = block_miss ? 1'h0 : T452;
  assign T452 = T459 ? 1'h0 : T453;
  assign T453 = T458 ? 1'h0 : T454;
  assign T454 = T455 == 1'h0;
  assign T455 = T457 & T456;
  assign T456 = io_cpu_req_bits_phys ^ 1'h1;
  assign T457 = dtlb_io_req_ready ^ 1'h1;
  assign T458 = metaReadArb_io_in_4_ready ^ 1'h1;
  assign T459 = readArb_io_in_3_ready ^ 1'h1;
  assign T460 = reset ? 1'h0 : T461;
  assign T461 = T462 & s2_nack_miss;
  assign T462 = s2_valid | block_miss;
  WritebackUnit wb(.clk(clk), .reset(reset),
       .io_req_ready( wb_io_req_ready ),
       .io_req_valid( wbArb_io_out_valid ),
       .io_req_bits_tag( wbArb_io_out_bits_tag ),
       .io_req_bits_idx( wbArb_io_out_bits_idx ),
       .io_req_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_req_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_req_bits_master_xact_id( wbArb_io_out_bits_master_xact_id ),
       .io_req_bits_r_type( wbArb_io_out_bits_r_type ),
       .io_meta_read_ready( metaReadArb_io_in_3_ready ),
       .io_meta_read_valid( wb_io_meta_read_valid ),
       .io_meta_read_bits_idx( wb_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( wb_io_meta_read_bits_tag ),
       .io_data_req_ready( readArb_io_in_2_ready ),
       .io_data_req_valid( wb_io_data_req_valid ),
       .io_data_req_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_data_req_bits_addr( wb_io_data_req_bits_addr ),
       .io_data_resp( s2_data_corrected ),
       .io_release_ready( releaseArb_io_in_0_ready ),
       .io_release_valid( wb_io_release_valid ),
       .io_release_bits_addr( wb_io_release_bits_addr ),
       .io_release_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_release_bits_master_xact_id( wb_io_release_bits_master_xact_id ),
       .io_release_bits_data( wb_io_release_bits_data ),
       .io_release_bits_r_type( wb_io_release_bits_r_type )
  );
  ProbeUnit prober(.clk(clk), .reset(reset),
       .io_req_ready( prober_io_req_ready ),
       .io_req_valid( T335 ),
       .io_req_bits_addr( probe_bits_addr ),
       .io_req_bits_master_xact_id( probe_bits_master_xact_id ),
       .io_req_bits_p_type( probe_bits_p_type ),
       //.io_req_bits_client_xact_id(  )
       .io_rep_ready( releaseArb_io_in_1_ready ),
       .io_rep_valid( prober_io_rep_valid ),
       .io_rep_bits_addr( prober_io_rep_bits_addr ),
       .io_rep_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_rep_bits_master_xact_id( prober_io_rep_bits_master_xact_id ),
       .io_rep_bits_data( prober_io_rep_bits_data ),
       .io_rep_bits_r_type( prober_io_rep_bits_r_type ),
       .io_meta_read_ready( metaReadArb_io_in_2_ready ),
       .io_meta_read_valid( prober_io_meta_read_valid ),
       .io_meta_read_bits_idx( prober_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( prober_io_meta_read_bits_tag ),
       .io_meta_write_ready( metaWriteArb_io_in_1_ready ),
       .io_meta_write_valid( prober_io_meta_write_valid ),
       .io_meta_write_bits_idx( prober_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_wb_req_ready( wbArb_io_in_0_ready ),
       .io_wb_req_valid( prober_io_wb_req_valid ),
       .io_wb_req_bits_tag( prober_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( prober_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( prober_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_way_en( s2_tag_match_way ),
       .io_mshr_rdy( mshrs_io_probe_rdy ),
       .io_line_state_state( s2_hit_state_state )
  );
  `ifndef SYNTHESIS
    assign prober.io_req_bits_client_xact_id = {1{$random}};
  `endif
  MSHRFile mshrs(.clk(clk), .reset(reset),
       .io_req_ready( mshrs_io_req_ready ),
       .io_req_valid( T312 ),
       .io_req_bits_kill( s2_req_kill ),
       .io_req_bits_typ( s2_req_typ ),
       .io_req_bits_phys( s2_req_phys ),
       .io_req_bits_addr( s2_req_addr ),
       .io_req_bits_data( s2_req_data ),
       .io_req_bits_tag( s2_req_tag ),
       .io_req_bits_cmd( s2_req_cmd ),
       .io_req_bits_tag_match( T77 ),
       .io_req_bits_old_meta_tag( T303 ),
       .io_req_bits_old_meta_coh_state( T295 ),
       .io_req_bits_way_en( T290 ),
       .io_secondary_miss( mshrs_io_secondary_miss ),
       .io_mem_req_ready( T289 ),
       .io_mem_req_valid( mshrs_io_mem_req_valid ),
       .io_mem_req_bits_addr( mshrs_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( mshrs_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_data( mshrs_io_mem_req_bits_data ),
       .io_mem_req_bits_a_type( mshrs_io_mem_req_bits_a_type ),
       .io_mem_req_bits_write_mask( mshrs_io_mem_req_bits_write_mask ),
       .io_mem_req_bits_subword_addr( mshrs_io_mem_req_bits_subword_addr ),
       .io_mem_req_bits_atomic_opcode( mshrs_io_mem_req_bits_atomic_opcode ),
       .io_mem_resp_way_en( mshrs_io_mem_resp_way_en ),
       .io_mem_resp_addr( mshrs_io_mem_resp_addr ),
       //.io_mem_resp_wmask(  )
       //.io_mem_resp_data(  )
       .io_meta_read_ready( metaReadArb_io_in_1_ready ),
       .io_meta_read_valid( mshrs_io_meta_read_valid ),
       .io_meta_read_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_meta_read_bits_tag(  )
       .io_meta_write_ready( metaWriteArb_io_in_0_ready ),
       .io_meta_write_valid( mshrs_io_meta_write_valid ),
       .io_meta_write_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( readArb_io_in_1_ready ),
       .io_replay_valid( mshrs_io_replay_valid ),
       .io_replay_bits_kill( mshrs_io_replay_bits_kill ),
       .io_replay_bits_typ( mshrs_io_replay_bits_typ ),
       .io_replay_bits_phys( mshrs_io_replay_bits_phys ),
       .io_replay_bits_addr( mshrs_io_replay_bits_addr ),
       .io_replay_bits_data( mshrs_io_replay_bits_data ),
       .io_replay_bits_tag( mshrs_io_replay_bits_tag ),
       .io_replay_bits_cmd( mshrs_io_replay_bits_cmd ),
       //.io_replay_bits_sdq_id(  )
       .io_mem_grant_valid( T288 ),
       .io_mem_grant_bits_header_src( FlowThroughSerializer_io_out_bits_header_src ),
       .io_mem_grant_bits_header_dst( FlowThroughSerializer_io_out_bits_header_dst ),
       .io_mem_grant_bits_payload_data( FlowThroughSerializer_io_out_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( FlowThroughSerializer_io_out_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( FlowThroughSerializer_io_out_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( FlowThroughSerializer_io_out_bits_payload_g_type ),
       .io_mem_finish_ready( io_mem_finish_ready ),
       .io_mem_finish_valid( mshrs_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( mshrs_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( mshrs_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( mshrs_io_mem_finish_bits_payload_master_xact_id ),
       .io_wb_req_ready( wbArb_io_in_1_ready ),
       .io_wb_req_valid( mshrs_io_wb_req_valid ),
       .io_wb_req_bits_tag( mshrs_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( mshrs_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( mshrs_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_probe_rdy( mshrs_io_probe_rdy ),
       .io_fence_rdy( mshrs_io_fence_rdy )
  );
  TLB dtlb(.clk(clk), .reset(reset),
       .io_req_ready( dtlb_io_req_ready ),
       .io_req_valid( T275 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T274 ),
       .io_req_bits_passthrough( s1_req_phys ),
       .io_req_bits_instruction( 1'h0 ),
       .io_resp_miss( dtlb_io_resp_miss ),
       //.io_resp_hit_idx(  )
       .io_resp_ppn( dtlb_io_resp_ppn ),
       .io_resp_xcpt_ld( dtlb_io_resp_xcpt_ld ),
       .io_resp_xcpt_st( dtlb_io_resp_xcpt_st ),
       //.io_resp_xcpt_if(  )
       .io_ptw_req_ready( io_cpu_ptw_req_ready ),
       .io_ptw_req_valid( dtlb_io_ptw_req_valid ),
       .io_ptw_req_bits( dtlb_io_ptw_req_bits ),
       .io_ptw_resp_valid( io_cpu_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_cpu_ptw_resp_bits_error ),
       .io_ptw_resp_bits_ppn( io_cpu_ptw_resp_bits_ppn ),
       .io_ptw_resp_bits_perm( io_cpu_ptw_resp_bits_perm ),
       .io_ptw_status_ip( io_cpu_ptw_status_ip ),
       .io_ptw_status_im( io_cpu_ptw_status_im ),
       .io_ptw_status_zero( io_cpu_ptw_status_zero ),
       .io_ptw_status_er( io_cpu_ptw_status_er ),
       .io_ptw_status_vm( io_cpu_ptw_status_vm ),
       .io_ptw_status_s64( io_cpu_ptw_status_s64 ),
       .io_ptw_status_u64( io_cpu_ptw_status_u64 ),
       .io_ptw_status_ef( io_cpu_ptw_status_ef ),
       .io_ptw_status_pei( io_cpu_ptw_status_pei ),
       .io_ptw_status_ei( io_cpu_ptw_status_ei ),
       .io_ptw_status_ps( io_cpu_ptw_status_ps ),
       .io_ptw_status_s( io_cpu_ptw_status_s ),
       .io_ptw_invalidate( io_cpu_ptw_invalidate ),
       .io_ptw_sret( io_cpu_ptw_sret )
  );
  MetadataArray meta(.clk(clk), .reset(reset),
       .io_read_ready( meta_io_read_ready ),
       .io_read_valid( metaReadArb_io_out_valid ),
       .io_read_bits_idx( metaReadArb_io_out_bits_idx ),
       .io_write_ready( meta_io_write_ready ),
       .io_write_valid( metaWriteArb_io_out_valid ),
       .io_write_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_write_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_write_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_write_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state ),
       .io_resp_0_tag( meta_io_resp_0_tag ),
       .io_resp_0_coh_state( meta_io_resp_0_coh_state )
  );
  Arbiter_7 metaReadArb(
       .io_in_4_ready( metaReadArb_io_in_4_ready ),
       .io_in_4_valid( io_cpu_req_valid ),
       .io_in_4_bits_idx( T266 ),
       .io_in_3_ready( metaReadArb_io_in_3_ready ),
       .io_in_3_valid( wb_io_meta_read_valid ),
       .io_in_3_bits_idx( wb_io_meta_read_bits_idx ),
       .io_in_2_ready( metaReadArb_io_in_2_ready ),
       .io_in_2_valid( prober_io_meta_read_valid ),
       .io_in_2_bits_idx( prober_io_meta_read_bits_idx ),
       .io_in_1_ready( metaReadArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_meta_read_valid ),
       .io_in_1_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_idx( T264 ),
       .io_out_ready( meta_io_read_ready ),
       .io_out_valid( metaReadArb_io_out_valid ),
       .io_out_bits_idx( metaReadArb_io_out_bits_idx )
       //.io_chosen(  )
  );
  Arbiter_1 metaWriteArb(
       .io_in_1_ready( metaWriteArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_meta_write_valid ),
       .io_in_1_bits_idx( prober_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( metaWriteArb_io_in_0_ready ),
       .io_in_0_valid( mshrs_io_meta_write_valid ),
       .io_in_0_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_out_ready( meta_io_write_ready ),
       .io_out_valid( metaWriteArb_io_out_valid ),
       .io_out_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_out_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_out_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  DataArray data(.clk(clk),
       //.io_read_ready(  )
       .io_read_valid( readArb_io_out_valid ),
       .io_read_bits_way_en( readArb_io_out_bits_way_en ),
       .io_read_bits_addr( readArb_io_out_bits_addr ),
       .io_write_ready( data_io_write_ready ),
       .io_write_valid( writeArb_io_out_valid ),
       .io_write_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_write_bits_addr( writeArb_io_out_bits_addr ),
       .io_write_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_write_bits_data( T260 ),
       .io_resp_0( data_io_resp_0 )
  );
  Arbiter_8 readArb(
       .io_in_3_ready( readArb_io_in_3_ready ),
       .io_in_3_valid( io_cpu_req_valid ),
       .io_in_3_bits_way_en( 1'h1 ),
       .io_in_3_bits_addr( T259 ),
       .io_in_2_ready( readArb_io_in_2_ready ),
       .io_in_2_valid( wb_io_data_req_valid ),
       .io_in_2_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_in_2_bits_addr( wb_io_data_req_bits_addr ),
       .io_in_1_ready( readArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_replay_valid ),
       .io_in_1_bits_way_en( 1'h1 ),
       .io_in_1_bits_addr( T258 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_way_en( 1'h1 ),
       .io_in_0_bits_addr( T257 ),
       .io_out_ready( T255 ),
       .io_out_valid( readArb_io_out_valid ),
       .io_out_bits_way_en( readArb_io_out_bits_way_en ),
       .io_out_bits_addr( readArb_io_out_bits_addr )
       //.io_chosen(  )
  );
  Arbiter_9 writeArb(
       .io_in_1_ready( writeArb_io_in_1_ready ),
       .io_in_1_valid( T251 ),
       .io_in_1_bits_way_en( mshrs_io_mem_resp_way_en ),
       .io_in_1_bits_addr( mshrs_io_mem_resp_addr ),
       .io_in_1_bits_wmask( 2'h3 ),
       .io_in_1_bits_data( T250 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s3_valid ),
       .io_in_0_bits_way_en( s3_way ),
       .io_in_0_bits_addr( T248 ),
       .io_in_0_bits_wmask( T245 ),
       .io_in_0_bits_data( T244 ),
       .io_out_ready( data_io_write_ready ),
       .io_out_valid( writeArb_io_out_valid ),
       .io_out_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_out_bits_addr( writeArb_io_out_bits_addr ),
       .io_out_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_out_bits_data( writeArb_io_out_bits_data )
       //.io_chosen(  )
  );
  AMOALU amoalu(
       .io_addr( T243 ),
       .io_cmd( T242 ),
       .io_typ( s2_req_typ ),
       .io_lhs( T103 ),
       .io_rhs( s2_req_data ),
       .io_out( amoalu_io_out )
  );
  Arbiter_10 releaseArb(
       .io_in_1_ready( releaseArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_rep_valid ),
       .io_in_1_bits_addr( prober_io_rep_bits_addr ),
       .io_in_1_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_in_1_bits_master_xact_id( prober_io_rep_bits_master_xact_id ),
       .io_in_1_bits_data( prober_io_rep_bits_data ),
       .io_in_1_bits_r_type( prober_io_rep_bits_r_type ),
       .io_in_0_ready( releaseArb_io_in_0_ready ),
       .io_in_0_valid( wb_io_release_valid ),
       .io_in_0_bits_addr( wb_io_release_bits_addr ),
       .io_in_0_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_in_0_bits_master_xact_id( wb_io_release_bits_master_xact_id ),
       .io_in_0_bits_data( wb_io_release_bits_data ),
       .io_in_0_bits_r_type( wb_io_release_bits_r_type ),
       .io_out_ready( T5 ),
       .io_out_valid( releaseArb_io_out_valid ),
       .io_out_bits_addr( releaseArb_io_out_bits_addr ),
       .io_out_bits_client_xact_id( releaseArb_io_out_bits_client_xact_id ),
       .io_out_bits_master_xact_id( releaseArb_io_out_bits_master_xact_id ),
       .io_out_bits_data( releaseArb_io_out_bits_data ),
       .io_out_bits_r_type( releaseArb_io_out_bits_r_type )
       //.io_chosen(  )
  );
  FlowThroughSerializer_1 FlowThroughSerializer(.clk(clk), .reset(reset),
       .io_in_ready( FlowThroughSerializer_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_header_src( io_mem_grant_bits_header_src ),
       .io_in_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_in_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_in_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_in_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_in_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_out_ready( T0 ),
       .io_out_valid( FlowThroughSerializer_io_out_valid ),
       .io_out_bits_header_src( FlowThroughSerializer_io_out_bits_header_src ),
       .io_out_bits_header_dst( FlowThroughSerializer_io_out_bits_header_dst ),
       .io_out_bits_payload_data( FlowThroughSerializer_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( FlowThroughSerializer_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( FlowThroughSerializer_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( FlowThroughSerializer_io_out_bits_payload_g_type )
       //.io_cnt(  )
       //.io_done(  )
  );
  Arbiter_4 wbArb(
       .io_in_1_ready( wbArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_wb_req_valid ),
       .io_in_1_bits_tag( mshrs_io_wb_req_bits_tag ),
       .io_in_1_bits_idx( mshrs_io_wb_req_bits_idx ),
       .io_in_1_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_in_1_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_master_xact_id( mshrs_io_wb_req_bits_master_xact_id ),
       .io_in_1_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_in_0_ready( wbArb_io_in_0_ready ),
       .io_in_0_valid( prober_io_wb_req_valid ),
       .io_in_0_bits_tag( prober_io_wb_req_bits_tag ),
       .io_in_0_bits_idx( prober_io_wb_req_bits_idx ),
       .io_in_0_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_in_0_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_master_xact_id( prober_io_wb_req_bits_master_xact_id ),
       .io_in_0_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_out_ready( wb_io_req_ready ),
       .io_out_valid( wbArb_io_out_valid ),
       .io_out_bits_tag( wbArb_io_out_bits_tag ),
       .io_out_bits_idx( wbArb_io_out_bits_idx ),
       .io_out_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_out_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_out_bits_master_xact_id( wbArb_io_out_bits_master_xact_id ),
       .io_out_bits_r_type( wbArb_io_out_bits_r_type )
       //.io_chosen(  )
  );

  always @(posedge clk) begin
    if(T101) begin
      s2_req_data <= s1_req_data;
    end else if(T11) begin
      s2_req_data <= T8;
    end
    if(reset) begin
      s1_replay <= 1'h0;
    end else begin
      s1_replay <= T10;
    end
    if(s2_recycle) begin
      s1_req_cmd <= s2_req_cmd;
    end else if(mshrs_io_replay_valid) begin
      s1_req_cmd <= mshrs_io_replay_bits_cmd;
    end else if(io_cpu_req_valid) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if(s1_clk_en) begin
      s2_req_cmd <= s1_req_cmd;
    end
    s1_clk_en <= metaReadArb_io_out_valid;
    if(reset) begin
      s2_recycle_next <= 1'h0;
    end else if(T93) begin
      s2_recycle_next <= T21;
    end
    if(s1_clk_en) begin
      s2_req_addr <= T29;
    end
    if(s2_recycle) begin
      s1_req_addr <= s2_req_addr;
    end else if(mshrs_io_replay_valid) begin
      s1_req_addr <= mshrs_io_replay_bits_addr;
    end else if(prober_io_meta_read_valid) begin
      s1_req_addr <= T39;
    end else if(wb_io_meta_read_valid) begin
      s1_req_addr <= T36;
    end else if(io_cpu_req_valid) begin
      s1_req_addr <= io_cpu_req_bits_addr;
    end
    if(s1_clk_en) begin
      s2_hit_state_state <= meta_io_resp_0_coh_state;
    end
    if(s1_clk_en) begin
      s2_tag_match_way <= s1_tag_match_way;
    end
    if(reset) begin
      R86 <= 1'h0;
    end else begin
      R86 <= s1_replay;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s1_valid_masked;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T91;
    end
    if(s2_recycle) begin
      s1_req_data <= s2_req_data;
    end else if(mshrs_io_replay_valid) begin
      s1_req_data <= mshrs_io_replay_bits_data;
    end else if(io_cpu_req_valid) begin
      s1_req_data <= io_cpu_req_bits_data;
    end
    if(s1_clk_en) begin
      s1_recycled <= s2_recycle;
    end
    R109 <= T110;
    if(T114) begin
      R116 <= T118;
    end
    if(T217) begin
      s2_store_bypass_data <= T122;
    end
    if(T142) begin
      s4_req_data <= s3_req_data;
    end
    s3_req_data <= T125;
    if(reset) begin
      s3_valid <= 1'h0;
    end else begin
      s3_valid <= T144;
    end
    if(T159) begin
      lrsc_addr <= T158;
    end
    if(T173) begin
      s2_nack_hit <= s1_nack;
    end
    if(reset) begin
      lrsc_count <= 5'h0;
    end else if(io_cpu_ptw_sret) begin
      lrsc_count <= 5'h0;
    end else if(T183) begin
      lrsc_count <= 5'h0;
    end else if(T181) begin
      lrsc_count <= 5'h1f;
    end else if(T174) begin
      lrsc_count <= T180;
    end
    if(T129) begin
      s3_req_cmd <= s2_req_cmd;
    end
    if(T129) begin
      s3_req_addr <= s2_req_addr;
    end
    if(T142) begin
      s4_req_cmd <= s3_req_cmd;
    end
    if(T142) begin
      s4_req_addr <= s3_req_addr;
    end
    if(reset) begin
      s4_valid <= 1'h0;
    end else begin
      s4_valid <= s3_valid;
    end
    if(T217) begin
      s2_store_bypass <= 1'h1;
    end else if(s1_clk_en) begin
      s2_store_bypass <= 1'h0;
    end
    if(s1_clk_en) begin
      s2_req_typ <= s1_req_typ;
    end
    if(s2_recycle) begin
      s1_req_typ <= s2_req_typ;
    end else if(mshrs_io_replay_valid) begin
      s1_req_typ <= mshrs_io_replay_bits_typ;
    end else if(io_cpu_req_valid) begin
      s1_req_typ <= io_cpu_req_bits_typ;
    end
    if(T129) begin
      s3_way <= s2_tag_match_way;
    end
    if(s2_recycle) begin
      s1_req_phys <= s2_req_phys;
    end else if(mshrs_io_replay_valid) begin
      s1_req_phys <= mshrs_io_replay_bits_phys;
    end else if(prober_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(wb_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s1_req_phys <= io_cpu_req_bits_phys;
    end
    if(s1_clk_en) begin
      s2_req_phys <= s1_req_phys;
    end
    if(s1_clk_en) begin
      R292 <= 1'h0;
    end
    if(s1_clk_en) begin
      s2_repl_meta_coh_state <= meta_io_resp_0_coh_state;
    end
    if(s1_clk_en) begin
      s2_repl_meta_tag <= meta_io_resp_0_tag;
    end
    if(s1_clk_en) begin
      s2_req_tag <= s1_req_tag;
    end
    if(s2_recycle) begin
      s1_req_tag <= s2_req_tag;
    end else if(mshrs_io_replay_valid) begin
      s1_req_tag <= mshrs_io_replay_bits_tag;
    end else if(io_cpu_req_valid) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if(s1_clk_en) begin
      s2_req_kill <= s1_req_kill;
    end
    if(s2_recycle) begin
      s1_req_kill <= s2_req_kill;
    end else if(mshrs_io_replay_valid) begin
      s1_req_kill <= mshrs_io_replay_bits_kill;
    end else if(io_cpu_req_valid) begin
      s1_req_kill <= io_cpu_req_bits_kill;
    end
    if(reset) begin
      block_miss <= 1'h0;
    end else begin
      block_miss <= T461;
    end
  end
endmodule

module RRArbiter_0(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [29:0] io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [29:0] io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output[29:0] io_out_bits,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  R5;
  wire T6;
  wire T7;
  wire T8;
  wire[29:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R5 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T3 ? 1'h1 : T2;
  assign T2 = io_in_0_valid == 1'h0;
  assign T3 = io_in_1_valid & T4;
  assign T4 = R5 < 1'h1;
  assign T6 = reset ? 1'h0 : T7;
  assign T7 = T8 ? T0 : R5;
  assign T8 = io_out_ready & io_out_valid;
  assign io_out_bits = T9;
  assign T9 = T10 ? io_in_1_bits : io_in_0_bits;
  assign T10 = T0;
  assign io_out_valid = T11;
  assign T11 = T10 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T12;
  assign T12 = T13 & io_out_ready;
  assign T13 = T14;
  assign T14 = T21 | T15;
  assign T15 = T16 ^ 1'h1;
  assign T16 = T19 | T17;
  assign T17 = io_in_1_valid & T18;
  assign T18 = R5 < 1'h1;
  assign T19 = io_in_0_valid & T20;
  assign T20 = R5 < 1'h0;
  assign T21 = R5 < 1'h0;
  assign io_in_1_ready = T22;
  assign T22 = T23 & io_out_ready;
  assign T23 = T24;
  assign T24 = T28 | T25;
  assign T25 = T26 ^ 1'h1;
  assign T26 = T27 | io_in_0_valid;
  assign T27 = T19 | T17;
  assign T28 = T30 & T29;
  assign T29 = R5 < 1'h1;
  assign T30 = T19 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R5 <= 1'h0;
    end else if(T8) begin
      R5 <= T0;
    end
  end
endmodule

module PTW(input clk, input reset,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input [29:0] io_requestor_1_req_bits,
    output io_requestor_1_resp_valid,
    output io_requestor_1_resp_bits_error,
    output[18:0] io_requestor_1_resp_bits_ppn,
    output[5:0] io_requestor_1_resp_bits_perm,
    output[7:0] io_requestor_1_status_ip,
    output[7:0] io_requestor_1_status_im,
    output[6:0] io_requestor_1_status_zero,
    output io_requestor_1_status_er,
    output io_requestor_1_status_vm,
    output io_requestor_1_status_s64,
    output io_requestor_1_status_u64,
    output io_requestor_1_status_ef,
    output io_requestor_1_status_pei,
    output io_requestor_1_status_ei,
    output io_requestor_1_status_ps,
    output io_requestor_1_status_s,
    output io_requestor_1_invalidate,
    output io_requestor_1_sret,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input [29:0] io_requestor_0_req_bits,
    output io_requestor_0_resp_valid,
    output io_requestor_0_resp_bits_error,
    output[18:0] io_requestor_0_resp_bits_ppn,
    output[5:0] io_requestor_0_resp_bits_perm,
    output[7:0] io_requestor_0_status_ip,
    output[7:0] io_requestor_0_status_im,
    output[6:0] io_requestor_0_status_zero,
    output io_requestor_0_status_er,
    output io_requestor_0_status_vm,
    output io_requestor_0_status_s64,
    output io_requestor_0_status_u64,
    output io_requestor_0_status_ef,
    output io_requestor_0_status_pei,
    output io_requestor_0_status_ei,
    output io_requestor_0_status_ps,
    output io_requestor_0_status_s,
    output io_requestor_0_invalidate,
    output io_requestor_0_sret,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output io_mem_req_bits_kill,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_phys,
    output[43:0] io_mem_req_bits_addr,
    //output[63:0] io_mem_req_bits_data
    //output[7:0] io_mem_req_bits_tag
    output[4:0] io_mem_req_bits_cmd,
    input  io_mem_resp_valid,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input [2:0] io_mem_resp_bits_typ,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data,
    input [63:0] io_mem_resp_bits_data_subword,
    input [7:0] io_mem_resp_bits_tag,
    input [3:0] io_mem_resp_bits_cmd,
    input [43:0] io_mem_resp_bits_addr,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [7:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_ptw_req_ready
    //input  io_mem_ptw_req_valid
    //input [29:0] io_mem_ptw_req_bits
    //output io_mem_ptw_resp_valid
    //output io_mem_ptw_resp_bits_error
    //output[18:0] io_mem_ptw_resp_bits_ppn
    //output[5:0] io_mem_ptw_resp_bits_perm
    //output[7:0] io_mem_ptw_status_ip
    //output[7:0] io_mem_ptw_status_im
    //output[6:0] io_mem_ptw_status_zero
    //output io_mem_ptw_status_er
    //output io_mem_ptw_status_vm
    //output io_mem_ptw_status_s64
    //output io_mem_ptw_status_u64
    //output io_mem_ptw_status_ef
    //output io_mem_ptw_status_pei
    //output io_mem_ptw_status_ei
    //output io_mem_ptw_status_ps
    //output io_mem_ptw_status_s
    //output io_mem_ptw_invalidate
    //output io_mem_ptw_sret
    input  io_mem_ordered,
    input [31:0] io_dpath_ptbr,
    input  io_dpath_invalidate,
    input  io_dpath_sret,
    input [7:0] io_dpath_status_ip,
    input [7:0] io_dpath_status_im,
    input [6:0] io_dpath_status_zero,
    input  io_dpath_status_er,
    input  io_dpath_status_vm,
    input  io_dpath_status_s64,
    input  io_dpath_status_u64,
    input  io_dpath_status_ef,
    input  io_dpath_status_pei,
    input  io_dpath_status_ei,
    input  io_dpath_status_ps,
    input  io_dpath_status_s
);

  wire T0;
  reg [2:0] state;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire T10;
  wire arb_io_out_valid;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  reg [1:0] count;
  wire[1:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire T29;
  wire T30;
  wire[43:0] T31;
  wire[31:0] T32;
  wire[28:0] T33;
  wire[28:0] T34;
  wire[9:0] T35;
  wire[9:0] T36;
  wire[9:0] T37;
  wire[9:0] T38;
  reg [29:0] r_req_vpn;
  wire[29:0] T39;
  wire[29:0] arb_io_out_bits;
  wire T40;
  wire[9:0] T41;
  wire[19:0] T42;
  wire T43;
  wire[1:0] T44;
  wire[9:0] T45;
  wire[29:0] T46;
  wire T47;
  wire[18:0] T48;
  reg [63:0] r_pte;
  wire[63:0] T49;
  wire[63:0] T50;
  wire[63:0] T51;
  wire[31:0] T52;
  wire[12:0] T53;
  wire[18:0] T54;
  wire T55;
  wire[5:0] T56;
  wire[18:0] T57;
  wire[30:0] T58;
  wire[30:0] T59;
  wire[30:0] T60;
  wire[30:0] T61;
  wire[19:0] T62;
  wire[10:0] T63;
  wire[30:0] r_resp_ppn;
  wire[30:0] T64;
  wire[9:0] T65;
  wire[20:0] T66;
  wire T67;
  wire[1:0] T68;
  wire T69;
  wire resp_err;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  reg  r_req_dest;
  wire T74;
  wire arb_io_chosen;
  wire resp_val;
  wire T75;
  wire T76;
  wire arb_io_in_0_ready;
  wire[5:0] T77;
  wire[18:0] T78;
  wire[30:0] T79;
  wire T80;
  wire T81;
  wire arb_io_in_1_ready;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    count = {1{$random}};
    r_req_vpn = {1{$random}};
    r_pte = {2{$random}};
    r_req_dest = {1{$random}};
  end
`endif

  assign T0 = state == 3'h0;
  assign T1 = reset ? 3'h0 : T2;
  assign T2 = T30 ? 3'h0 : T3;
  assign T3 = T29 ? 3'h0 : T4;
  assign T4 = T22 ? 3'h1 : T5;
  assign T5 = T17 ? 3'h3 : T6;
  assign T6 = T16 ? 3'h4 : T7;
  assign T7 = T14 ? 3'h1 : T8;
  assign T8 = T12 ? 3'h2 : T9;
  assign T9 = T10 ? 3'h1 : state;
  assign T10 = T11 & arb_io_out_valid;
  assign T11 = 3'h0 == state;
  assign T12 = T13 & io_mem_req_ready;
  assign T13 = 3'h1 == state;
  assign T14 = T15 & io_mem_resp_bits_nack;
  assign T15 = 3'h2 == state;
  assign T16 = T15 & io_mem_resp_valid;
  assign T17 = T20 & T18;
  assign T18 = T19 ^ 1'h1;
  assign T19 = io_mem_resp_bits_data[1'h1:1'h1];
  assign T20 = T16 & T21;
  assign T21 = io_mem_resp_bits_data[1'h0:1'h0];
  assign T22 = T20 & T23;
  assign T23 = T28 & T24;
  assign T24 = count < 2'h2;
  assign T25 = T22 ? T27 : T26;
  assign T26 = T11 ? 2'h0 : count;
  assign T27 = count + 2'h1;
  assign T28 = T18 ^ 1'h1;
  assign T29 = 3'h3 == state;
  assign T30 = 3'h4 == state;
  assign io_mem_req_bits_cmd = 5'h0;
  assign io_mem_req_bits_addr = T31;
  assign T31 = {12'h0, T32};
  assign T32 = T33 << 2'h3;
  assign T33 = T34;
  assign T34 = {T48, T35};
  assign T35 = T47 ? T45 : T36;
  assign T36 = T43 ? T41 : T37;
  assign T37 = T38[4'h9:1'h0];
  assign T38 = r_req_vpn >> 5'h14;
  assign T39 = T40 ? arb_io_out_bits : r_req_vpn;
  assign T40 = T0 & arb_io_out_valid;
  assign T41 = T42[4'h9:1'h0];
  assign T42 = r_req_vpn >> 4'ha;
  assign T43 = T44[1'h0:1'h0];
  assign T44 = count;
  assign T45 = T46[4'h9:1'h0];
  assign T46 = r_req_vpn >> 1'h0;
  assign T47 = T44[1'h1:1'h1];
  assign T48 = r_pte[5'h1f:4'hd];
  assign T49 = io_mem_resp_valid ? io_mem_resp_bits_data : T50;
  assign T50 = T40 ? T51 : r_pte;
  assign T51 = {32'h0, T52};
  assign T52 = {T54, T53};
  assign T53 = io_mem_resp_bits_data[4'hc:1'h0];
  assign T54 = io_dpath_ptbr[5'h1f:4'hd];
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_bits_typ = 3'h3;
  assign io_mem_req_bits_kill = 1'h0;
  assign io_mem_req_valid = T55;
  assign T55 = state == 3'h1;
  assign io_requestor_0_sret = io_dpath_sret;
  assign io_requestor_0_invalidate = io_dpath_invalidate;
  assign io_requestor_0_status_s = io_dpath_status_s;
  assign io_requestor_0_status_ps = io_dpath_status_ps;
  assign io_requestor_0_status_ei = io_dpath_status_ei;
  assign io_requestor_0_status_pei = io_dpath_status_pei;
  assign io_requestor_0_status_ef = io_dpath_status_ef;
  assign io_requestor_0_status_u64 = io_dpath_status_u64;
  assign io_requestor_0_status_s64 = io_dpath_status_s64;
  assign io_requestor_0_status_vm = io_dpath_status_vm;
  assign io_requestor_0_status_er = io_dpath_status_er;
  assign io_requestor_0_status_zero = io_dpath_status_zero;
  assign io_requestor_0_status_im = io_dpath_status_im;
  assign io_requestor_0_status_ip = io_dpath_status_ip;
  assign io_requestor_0_resp_bits_perm = T56;
  assign T56 = r_pte[4'h8:2'h3];
  assign io_requestor_0_resp_bits_ppn = T57;
  assign T57 = T58[5'h12:1'h0];
  assign T58 = T59;
  assign T59 = T69 ? r_resp_ppn : T60;
  assign T60 = T67 ? T64 : T61;
  assign T61 = {T63, T62};
  assign T62 = r_req_vpn[5'h13:1'h0];
  assign T63 = r_resp_ppn >> 5'h14;
  assign r_resp_ppn = io_mem_req_bits_addr >> 4'hd;
  assign T64 = {T66, T65};
  assign T65 = r_req_vpn[4'h9:1'h0];
  assign T66 = r_resp_ppn >> 4'ha;
  assign T67 = T68[1'h0:1'h0];
  assign T68 = count;
  assign T69 = T68[1'h1:1'h1];
  assign io_requestor_0_resp_bits_error = resp_err;
  assign resp_err = T71 | T70;
  assign T70 = state == 3'h2;
  assign T71 = state == 3'h4;
  assign io_requestor_0_resp_valid = T72;
  assign T72 = resp_val & T73;
  assign T73 = r_req_dest == 1'h0;
  assign T74 = T40 ? arb_io_chosen : r_req_dest;
  assign resp_val = T76 | T75;
  assign T75 = state == 3'h4;
  assign T76 = state == 3'h3;
  assign io_requestor_0_req_ready = arb_io_in_0_ready;
  assign io_requestor_1_sret = io_dpath_sret;
  assign io_requestor_1_invalidate = io_dpath_invalidate;
  assign io_requestor_1_status_s = io_dpath_status_s;
  assign io_requestor_1_status_ps = io_dpath_status_ps;
  assign io_requestor_1_status_ei = io_dpath_status_ei;
  assign io_requestor_1_status_pei = io_dpath_status_pei;
  assign io_requestor_1_status_ef = io_dpath_status_ef;
  assign io_requestor_1_status_u64 = io_dpath_status_u64;
  assign io_requestor_1_status_s64 = io_dpath_status_s64;
  assign io_requestor_1_status_vm = io_dpath_status_vm;
  assign io_requestor_1_status_er = io_dpath_status_er;
  assign io_requestor_1_status_zero = io_dpath_status_zero;
  assign io_requestor_1_status_im = io_dpath_status_im;
  assign io_requestor_1_status_ip = io_dpath_status_ip;
  assign io_requestor_1_resp_bits_perm = T77;
  assign T77 = r_pte[4'h8:2'h3];
  assign io_requestor_1_resp_bits_ppn = T78;
  assign T78 = T79[5'h12:1'h0];
  assign T79 = T59;
  assign io_requestor_1_resp_bits_error = resp_err;
  assign io_requestor_1_resp_valid = T80;
  assign T80 = resp_val & T81;
  assign T81 = r_req_dest == 1'h1;
  assign io_requestor_1_req_ready = arb_io_in_1_ready;
  RRArbiter_0 arb(.clk(clk), .reset(reset),
       .io_in_1_ready( arb_io_in_1_ready ),
       .io_in_1_valid( io_requestor_1_req_valid ),
       .io_in_1_bits( io_requestor_1_req_bits ),
       .io_in_0_ready( arb_io_in_0_ready ),
       .io_in_0_valid( io_requestor_0_req_valid ),
       .io_in_0_bits( io_requestor_0_req_bits ),
       .io_out_ready( T0 ),
       .io_out_valid( arb_io_out_valid ),
       .io_out_bits( arb_io_out_bits ),
       .io_chosen( arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T30) begin
      state <= 3'h0;
    end else if(T29) begin
      state <= 3'h0;
    end else if(T22) begin
      state <= 3'h1;
    end else if(T17) begin
      state <= 3'h3;
    end else if(T16) begin
      state <= 3'h4;
    end else if(T14) begin
      state <= 3'h1;
    end else if(T12) begin
      state <= 3'h2;
    end else if(T10) begin
      state <= 3'h1;
    end
    if(T22) begin
      count <= T27;
    end else if(T11) begin
      count <= 2'h0;
    end
    if(T40) begin
      r_req_vpn <= arb_io_out_bits;
    end
    if(io_mem_resp_valid) begin
      r_pte <= io_mem_resp_bits_data;
    end else if(T40) begin
      r_pte <= T51;
    end
    if(T40) begin
      r_req_dest <= arb_io_chosen;
    end
  end
endmodule

module HellaCacheArbiter(input clk,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input  io_requestor_1_req_bits_kill,
    input [2:0] io_requestor_1_req_bits_typ,
    input  io_requestor_1_req_bits_phys,
    input [43:0] io_requestor_1_req_bits_addr,
    input [63:0] io_requestor_1_req_bits_data,
    input [7:0] io_requestor_1_req_bits_tag,
    input [4:0] io_requestor_1_req_bits_cmd,
    output io_requestor_1_resp_valid,
    output io_requestor_1_resp_bits_nack,
    output io_requestor_1_resp_bits_replay,
    output[2:0] io_requestor_1_resp_bits_typ,
    output io_requestor_1_resp_bits_has_data,
    output[63:0] io_requestor_1_resp_bits_data,
    output[63:0] io_requestor_1_resp_bits_data_subword,
    output[7:0] io_requestor_1_resp_bits_tag,
    output[3:0] io_requestor_1_resp_bits_cmd,
    output[43:0] io_requestor_1_resp_bits_addr,
    output[63:0] io_requestor_1_resp_bits_store_data,
    output io_requestor_1_replay_next_valid,
    output[7:0] io_requestor_1_replay_next_bits,
    output io_requestor_1_xcpt_ma_ld,
    output io_requestor_1_xcpt_ma_st,
    output io_requestor_1_xcpt_pf_ld,
    output io_requestor_1_xcpt_pf_st,
    //input  io_requestor_1_ptw_req_ready
    //output io_requestor_1_ptw_req_valid
    //output[29:0] io_requestor_1_ptw_req_bits
    //input  io_requestor_1_ptw_resp_valid
    //input  io_requestor_1_ptw_resp_bits_error
    //input [18:0] io_requestor_1_ptw_resp_bits_ppn
    //input [5:0] io_requestor_1_ptw_resp_bits_perm
    //input [7:0] io_requestor_1_ptw_status_ip
    //input [7:0] io_requestor_1_ptw_status_im
    //input [6:0] io_requestor_1_ptw_status_zero
    //input  io_requestor_1_ptw_status_er
    //input  io_requestor_1_ptw_status_vm
    //input  io_requestor_1_ptw_status_s64
    //input  io_requestor_1_ptw_status_u64
    //input  io_requestor_1_ptw_status_ef
    //input  io_requestor_1_ptw_status_pei
    //input  io_requestor_1_ptw_status_ei
    //input  io_requestor_1_ptw_status_ps
    //input  io_requestor_1_ptw_status_s
    //input  io_requestor_1_ptw_invalidate
    //input  io_requestor_1_ptw_sret
    output io_requestor_1_ordered,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input  io_requestor_0_req_bits_kill,
    input [2:0] io_requestor_0_req_bits_typ,
    input  io_requestor_0_req_bits_phys,
    input [43:0] io_requestor_0_req_bits_addr,
    input [63:0] io_requestor_0_req_bits_data,
    input [7:0] io_requestor_0_req_bits_tag,
    input [4:0] io_requestor_0_req_bits_cmd,
    output io_requestor_0_resp_valid,
    output io_requestor_0_resp_bits_nack,
    output io_requestor_0_resp_bits_replay,
    output[2:0] io_requestor_0_resp_bits_typ,
    output io_requestor_0_resp_bits_has_data,
    output[63:0] io_requestor_0_resp_bits_data,
    output[63:0] io_requestor_0_resp_bits_data_subword,
    output[7:0] io_requestor_0_resp_bits_tag,
    output[3:0] io_requestor_0_resp_bits_cmd,
    output[43:0] io_requestor_0_resp_bits_addr,
    output[63:0] io_requestor_0_resp_bits_store_data,
    output io_requestor_0_replay_next_valid,
    output[7:0] io_requestor_0_replay_next_bits,
    output io_requestor_0_xcpt_ma_ld,
    output io_requestor_0_xcpt_ma_st,
    output io_requestor_0_xcpt_pf_ld,
    output io_requestor_0_xcpt_pf_st,
    //input  io_requestor_0_ptw_req_ready
    //output io_requestor_0_ptw_req_valid
    //output[29:0] io_requestor_0_ptw_req_bits
    //input  io_requestor_0_ptw_resp_valid
    //input  io_requestor_0_ptw_resp_bits_error
    //input [18:0] io_requestor_0_ptw_resp_bits_ppn
    //input [5:0] io_requestor_0_ptw_resp_bits_perm
    //input [7:0] io_requestor_0_ptw_status_ip
    //input [7:0] io_requestor_0_ptw_status_im
    //input [6:0] io_requestor_0_ptw_status_zero
    //input  io_requestor_0_ptw_status_er
    //input  io_requestor_0_ptw_status_vm
    //input  io_requestor_0_ptw_status_s64
    //input  io_requestor_0_ptw_status_u64
    //input  io_requestor_0_ptw_status_ef
    //input  io_requestor_0_ptw_status_pei
    //input  io_requestor_0_ptw_status_ei
    //input  io_requestor_0_ptw_status_ps
    //input  io_requestor_0_ptw_status_s
    //input  io_requestor_0_ptw_invalidate
    //input  io_requestor_0_ptw_sret
    output io_requestor_0_ordered,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output io_mem_req_bits_kill,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_phys,
    output[43:0] io_mem_req_bits_addr,
    output[63:0] io_mem_req_bits_data,
    output[7:0] io_mem_req_bits_tag,
    output[4:0] io_mem_req_bits_cmd,
    input  io_mem_resp_valid,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input [2:0] io_mem_resp_bits_typ,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data,
    input [63:0] io_mem_resp_bits_data_subword,
    input [7:0] io_mem_resp_bits_tag,
    input [3:0] io_mem_resp_bits_cmd,
    input [43:0] io_mem_resp_bits_addr,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [7:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_ptw_req_ready
    input  io_mem_ptw_req_valid,
    input [29:0] io_mem_ptw_req_bits,
    //output io_mem_ptw_resp_valid
    //output io_mem_ptw_resp_bits_error
    //output[18:0] io_mem_ptw_resp_bits_ppn
    //output[5:0] io_mem_ptw_resp_bits_perm
    //output[7:0] io_mem_ptw_status_ip
    //output[7:0] io_mem_ptw_status_im
    //output[6:0] io_mem_ptw_status_zero
    //output io_mem_ptw_status_er
    //output io_mem_ptw_status_vm
    //output io_mem_ptw_status_s64
    //output io_mem_ptw_status_u64
    //output io_mem_ptw_status_ef
    //output io_mem_ptw_status_pei
    //output io_mem_ptw_status_ei
    //output io_mem_ptw_status_ps
    //output io_mem_ptw_status_s
    //output io_mem_ptw_invalidate
    //output io_mem_ptw_sret
    input  io_mem_ordered
);

  wire[4:0] T0;
  wire[7:0] T1;
  wire[8:0] T2;
  wire[8:0] T3;
  wire[8:0] T4;
  wire[63:0] T5;
  reg  r_valid_0;
  wire[43:0] T6;
  wire T7;
  wire[2:0] T8;
  wire T9;
  wire T10;
  wire[7:0] T11;
  wire[6:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire[7:0] T16;
  wire[6:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire[7:0] T23;
  wire[6:0] T24;
  wire T25;
  wire T26;
  wire T27;
  wire[7:0] T28;
  wire[6:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    r_valid_0 = {1{$random}};
  end
`endif

  assign io_mem_req_bits_cmd = T0;
  assign T0 = io_requestor_0_req_valid ? io_requestor_0_req_bits_cmd : io_requestor_1_req_bits_cmd;
  assign io_mem_req_bits_tag = T1;
  assign T1 = T2[3'h7:1'h0];
  assign T2 = io_requestor_0_req_valid ? T4 : T3;
  assign T3 = {io_requestor_1_req_bits_tag, 1'h1};
  assign T4 = {io_requestor_0_req_bits_tag, 1'h0};
  assign io_mem_req_bits_data = T5;
  assign T5 = r_valid_0 ? io_requestor_0_req_bits_data : io_requestor_1_req_bits_data;
  assign io_mem_req_bits_addr = T6;
  assign T6 = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr;
  assign io_mem_req_bits_phys = T7;
  assign T7 = io_requestor_0_req_valid ? io_requestor_0_req_bits_phys : io_requestor_1_req_bits_phys;
  assign io_mem_req_bits_typ = T8;
  assign T8 = io_requestor_0_req_valid ? io_requestor_0_req_bits_typ : io_requestor_1_req_bits_typ;
  assign io_mem_req_bits_kill = T9;
  assign T9 = r_valid_0 ? io_requestor_0_req_bits_kill : io_requestor_1_req_bits_kill;
  assign io_mem_req_valid = T10;
  assign T10 = io_requestor_0_req_valid | io_requestor_1_req_valid;
  assign io_requestor_0_ordered = io_mem_ordered;
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_replay_next_bits = T11;
  assign T11 = {1'h0, T12};
  assign T12 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_0_replay_next_valid = T13;
  assign T13 = io_mem_replay_next_valid & T14;
  assign T14 = T15 == 1'h0;
  assign T15 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_0_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_0_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_0_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_0_resp_bits_tag = T16;
  assign T16 = {1'h0, T17};
  assign T17 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_0_resp_bits_data_subword = io_mem_resp_bits_data_subword;
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_0_resp_bits_replay = T18;
  assign T18 = io_mem_resp_bits_replay & T19;
  assign T19 = T20 == 1'h0;
  assign T20 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_0_resp_bits_nack = T21;
  assign T21 = io_mem_resp_bits_nack & T19;
  assign io_requestor_0_resp_valid = T22;
  assign T22 = io_mem_resp_valid & T19;
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_1_ordered = io_mem_ordered;
  assign io_requestor_1_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_1_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_1_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_1_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_1_replay_next_bits = T23;
  assign T23 = {1'h0, T24};
  assign T24 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_1_replay_next_valid = T25;
  assign T25 = io_mem_replay_next_valid & T26;
  assign T26 = T27 == 1'h1;
  assign T27 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_1_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_1_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_1_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_1_resp_bits_tag = T28;
  assign T28 = {1'h0, T29};
  assign T29 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_1_resp_bits_data_subword = io_mem_resp_bits_data_subword;
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_1_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_1_resp_bits_replay = T30;
  assign T30 = io_mem_resp_bits_replay & T31;
  assign T31 = T32 == 1'h1;
  assign T32 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_1_resp_bits_nack = T33;
  assign T33 = io_mem_resp_bits_nack & T31;
  assign io_requestor_1_resp_valid = T34;
  assign T34 = io_mem_resp_valid & T31;
  assign io_requestor_1_req_ready = T35;
  assign T35 = io_requestor_0_req_ready & T36;
  assign T36 = io_requestor_0_req_valid ^ 1'h1;

  always @(posedge clk) begin
    r_valid_0 <= io_requestor_0_req_valid;
  end
endmodule

module RRArbiter_1(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [3:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [3:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[3:0] io_out_bits_payload_client_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_a_type,
    output[5:0] io_out_bits_payload_write_mask,
    output[2:0] io_out_bits_payload_subword_addr,
    output[3:0] io_out_bits_payload_atomic_opcode,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  R5;
  wire T6;
  wire T7;
  wire T8;
  wire[3:0] T9;
  wire T10;
  wire[2:0] T11;
  wire[5:0] T12;
  wire[2:0] T13;
  wire[511:0] T14;
  wire[3:0] T15;
  wire[25:0] T16;
  wire[1:0] T17;
  wire[1:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R5 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T3 ? 1'h1 : T2;
  assign T2 = io_in_0_valid == 1'h0;
  assign T3 = io_in_1_valid & T4;
  assign T4 = R5 < 1'h1;
  assign T6 = reset ? 1'h0 : T7;
  assign T7 = T8 ? T0 : R5;
  assign T8 = io_out_ready & io_out_valid;
  assign io_out_bits_payload_atomic_opcode = T9;
  assign T9 = T10 ? io_in_1_bits_payload_atomic_opcode : io_in_0_bits_payload_atomic_opcode;
  assign T10 = T0;
  assign io_out_bits_payload_subword_addr = T11;
  assign T11 = T10 ? io_in_1_bits_payload_subword_addr : io_in_0_bits_payload_subword_addr;
  assign io_out_bits_payload_write_mask = T12;
  assign T12 = T10 ? io_in_1_bits_payload_write_mask : io_in_0_bits_payload_write_mask;
  assign io_out_bits_payload_a_type = T13;
  assign T13 = T10 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign io_out_bits_payload_data = T14;
  assign T14 = T10 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign io_out_bits_payload_client_xact_id = T15;
  assign T15 = T10 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign io_out_bits_payload_addr = T16;
  assign T16 = T10 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign io_out_bits_header_dst = T17;
  assign T17 = T10 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T18;
  assign T18 = T10 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T19;
  assign T19 = T10 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T20;
  assign T20 = T21 & io_out_ready;
  assign T21 = T22;
  assign T22 = T29 | T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = T27 | T25;
  assign T25 = io_in_1_valid & T26;
  assign T26 = R5 < 1'h1;
  assign T27 = io_in_0_valid & T28;
  assign T28 = R5 < 1'h0;
  assign T29 = R5 < 1'h0;
  assign io_in_1_ready = T30;
  assign T30 = T31 & io_out_ready;
  assign T31 = T32;
  assign T32 = T36 | T33;
  assign T33 = T34 ^ 1'h1;
  assign T34 = T35 | io_in_0_valid;
  assign T35 = T27 | T25;
  assign T36 = T38 & T37;
  assign T37 = R5 < 1'h1;
  assign T38 = T27 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R5 <= 1'h0;
    end else if(T8) begin
      R5 <= T0;
    end
  end
endmodule

module RRArbiter_2(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [3:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [3:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[3:0] io_out_bits_payload_master_xact_id,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  R5;
  wire T6;
  wire T7;
  wire T8;
  wire[3:0] T9;
  wire T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R5 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T3 ? 1'h1 : T2;
  assign T2 = io_in_0_valid == 1'h0;
  assign T3 = io_in_1_valid & T4;
  assign T4 = R5 < 1'h1;
  assign T6 = reset ? 1'h0 : T7;
  assign T7 = T8 ? T0 : R5;
  assign T8 = io_out_ready & io_out_valid;
  assign io_out_bits_payload_master_xact_id = T9;
  assign T9 = T10 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T10 = T0;
  assign io_out_bits_header_dst = T11;
  assign T11 = T10 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T12;
  assign T12 = T10 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T13;
  assign T13 = T10 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T14;
  assign T14 = T15 & io_out_ready;
  assign T15 = T16;
  assign T16 = T23 | T17;
  assign T17 = T18 ^ 1'h1;
  assign T18 = T21 | T19;
  assign T19 = io_in_1_valid & T20;
  assign T20 = R5 < 1'h1;
  assign T21 = io_in_0_valid & T22;
  assign T22 = R5 < 1'h0;
  assign T23 = R5 < 1'h0;
  assign io_in_1_ready = T24;
  assign T24 = T25 & io_out_ready;
  assign T25 = T26;
  assign T26 = T30 | T27;
  assign T27 = T28 ^ 1'h1;
  assign T28 = T29 | io_in_0_valid;
  assign T29 = T21 | T19;
  assign T30 = T32 & T31;
  assign T31 = R5 < 1'h1;
  assign T32 = T21 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R5 <= 1'h0;
    end else if(T8) begin
      R5 <= T0;
    end
  end
endmodule

module UncachedTileLinkIOArbiterThatAppendsArbiterId(input clk, input reset,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [1:0] io_in_1_acquire_bits_header_src,
    input [1:0] io_in_1_acquire_bits_header_dst,
    input [25:0] io_in_1_acquire_bits_payload_addr,
    input [3:0] io_in_1_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_1_acquire_bits_payload_data,
    input [2:0] io_in_1_acquire_bits_payload_a_type,
    input [5:0] io_in_1_acquire_bits_payload_write_mask,
    input [2:0] io_in_1_acquire_bits_payload_subword_addr,
    input [3:0] io_in_1_acquire_bits_payload_atomic_opcode,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_header_src,
    output[1:0] io_in_1_grant_bits_header_dst,
    output[511:0] io_in_1_grant_bits_payload_data,
    output[3:0] io_in_1_grant_bits_payload_client_xact_id,
    output[3:0] io_in_1_grant_bits_payload_master_xact_id,
    output[3:0] io_in_1_grant_bits_payload_g_type,
    output io_in_1_finish_ready,
    input  io_in_1_finish_valid,
    input [1:0] io_in_1_finish_bits_header_src,
    input [1:0] io_in_1_finish_bits_header_dst,
    input [3:0] io_in_1_finish_bits_payload_master_xact_id,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [1:0] io_in_0_acquire_bits_header_src,
    input [1:0] io_in_0_acquire_bits_header_dst,
    input [25:0] io_in_0_acquire_bits_payload_addr,
    input [3:0] io_in_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_0_acquire_bits_payload_data,
    input [2:0] io_in_0_acquire_bits_payload_a_type,
    input [5:0] io_in_0_acquire_bits_payload_write_mask,
    input [2:0] io_in_0_acquire_bits_payload_subword_addr,
    input [3:0] io_in_0_acquire_bits_payload_atomic_opcode,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_header_src,
    output[1:0] io_in_0_grant_bits_header_dst,
    output[511:0] io_in_0_grant_bits_payload_data,
    output[3:0] io_in_0_grant_bits_payload_client_xact_id,
    output[3:0] io_in_0_grant_bits_payload_master_xact_id,
    output[3:0] io_in_0_grant_bits_payload_g_type,
    output io_in_0_finish_ready,
    input  io_in_0_finish_valid,
    input [1:0] io_in_0_finish_bits_header_src,
    input [1:0] io_in_0_finish_bits_header_dst,
    input [3:0] io_in_0_finish_bits_payload_master_xact_id,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[1:0] io_out_acquire_bits_header_src,
    output[1:0] io_out_acquire_bits_header_dst,
    output[25:0] io_out_acquire_bits_payload_addr,
    output[3:0] io_out_acquire_bits_payload_client_xact_id,
    output[511:0] io_out_acquire_bits_payload_data,
    output[2:0] io_out_acquire_bits_payload_a_type,
    output[5:0] io_out_acquire_bits_payload_write_mask,
    output[2:0] io_out_acquire_bits_payload_subword_addr,
    output[3:0] io_out_acquire_bits_payload_atomic_opcode,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_header_src,
    input [1:0] io_out_grant_bits_header_dst,
    input [511:0] io_out_grant_bits_payload_data,
    input [3:0] io_out_grant_bits_payload_client_xact_id,
    input [3:0] io_out_grant_bits_payload_master_xact_id,
    input [3:0] io_out_grant_bits_payload_g_type,
    input  io_out_finish_ready,
    output io_out_finish_valid,
    output[1:0] io_out_finish_bits_header_src,
    output[1:0] io_out_finish_bits_header_dst,
    output[3:0] io_out_finish_bits_payload_master_xact_id
);

  wire[3:0] T0;
  wire[4:0] T1;
  wire[3:0] T2;
  wire[4:0] T3;
  wire[3:0] RRArbiter_1_io_out_bits_payload_master_xact_id;
  wire[1:0] RRArbiter_1_io_out_bits_header_dst;
  wire[1:0] RRArbiter_1_io_out_bits_header_src;
  wire RRArbiter_1_io_out_valid;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[3:0] RRArbiter_0_io_out_bits_payload_atomic_opcode;
  wire[2:0] RRArbiter_0_io_out_bits_payload_subword_addr;
  wire[5:0] RRArbiter_0_io_out_bits_payload_write_mask;
  wire[2:0] RRArbiter_0_io_out_bits_payload_a_type;
  wire[511:0] RRArbiter_0_io_out_bits_payload_data;
  wire[3:0] RRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[25:0] RRArbiter_0_io_out_bits_payload_addr;
  wire[1:0] RRArbiter_0_io_out_bits_header_dst;
  wire[1:0] RRArbiter_0_io_out_bits_header_src;
  wire RRArbiter_0_io_out_valid;
  wire RRArbiter_1_io_in_0_ready;
  wire[3:0] T12;
  wire[2:0] T13;
  wire T14;
  wire RRArbiter_0_io_in_0_ready;
  wire RRArbiter_1_io_in_1_ready;
  wire[3:0] T15;
  wire[2:0] T16;
  wire T17;
  wire RRArbiter_0_io_in_1_ready;


  assign T0 = T1[2'h3:1'h0];
  assign T1 = {io_in_0_acquire_bits_payload_client_xact_id, 1'h0};
  assign T2 = T3[2'h3:1'h0];
  assign T3 = {io_in_1_acquire_bits_payload_client_xact_id, 1'h1};
  assign io_out_finish_bits_payload_master_xact_id = RRArbiter_1_io_out_bits_payload_master_xact_id;
  assign io_out_finish_bits_header_dst = RRArbiter_1_io_out_bits_header_dst;
  assign io_out_finish_bits_header_src = RRArbiter_1_io_out_bits_header_src;
  assign io_out_finish_valid = RRArbiter_1_io_out_valid;
  assign io_out_grant_ready = T4;
  assign T4 = T9 ? io_in_1_grant_ready : T5;
  assign T5 = T6 ? io_in_0_grant_ready : 1'h0;
  assign T6 = T7 == 1'h0;
  assign T7 = T8;
  assign T8 = io_out_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign T9 = T10 == 1'h1;
  assign T10 = T11;
  assign T11 = io_out_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign io_out_acquire_bits_payload_atomic_opcode = RRArbiter_0_io_out_bits_payload_atomic_opcode;
  assign io_out_acquire_bits_payload_subword_addr = RRArbiter_0_io_out_bits_payload_subword_addr;
  assign io_out_acquire_bits_payload_write_mask = RRArbiter_0_io_out_bits_payload_write_mask;
  assign io_out_acquire_bits_payload_a_type = RRArbiter_0_io_out_bits_payload_a_type;
  assign io_out_acquire_bits_payload_data = RRArbiter_0_io_out_bits_payload_data;
  assign io_out_acquire_bits_payload_client_xact_id = RRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_acquire_bits_payload_addr = RRArbiter_0_io_out_bits_payload_addr;
  assign io_out_acquire_bits_header_dst = RRArbiter_0_io_out_bits_header_dst;
  assign io_out_acquire_bits_header_src = RRArbiter_0_io_out_bits_header_src;
  assign io_out_acquire_valid = RRArbiter_0_io_out_valid;
  assign io_in_0_finish_ready = RRArbiter_1_io_in_0_ready;
  assign io_in_0_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_0_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_0_grant_bits_payload_client_xact_id = T12;
  assign T12 = {1'h0, T13};
  assign T13 = io_out_grant_bits_payload_client_xact_id >> 1'h1;
  assign io_in_0_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_0_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_0_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_0_grant_valid = T14;
  assign T14 = T6 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = RRArbiter_0_io_in_0_ready;
  assign io_in_1_finish_ready = RRArbiter_1_io_in_1_ready;
  assign io_in_1_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_1_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_1_grant_bits_payload_client_xact_id = T15;
  assign T15 = {1'h0, T16};
  assign T16 = io_out_grant_bits_payload_client_xact_id >> 1'h1;
  assign io_in_1_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_1_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_1_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_1_grant_valid = T17;
  assign T17 = T9 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = RRArbiter_0_io_in_1_ready;
  RRArbiter_1 RRArbiter_0(.clk(clk), .reset(reset),
       .io_in_1_ready( RRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_header_src( io_in_1_acquire_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_acquire_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_acquire_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( T2 ),
       .io_in_1_bits_payload_data( io_in_1_acquire_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_acquire_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_acquire_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_acquire_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_acquire_bits_payload_atomic_opcode ),
       .io_in_0_ready( RRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_header_src( io_in_0_acquire_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_acquire_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_acquire_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( T0 ),
       .io_in_0_bits_payload_data( io_in_0_acquire_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_acquire_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_acquire_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_acquire_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_acquire_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( RRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( RRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( RRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( RRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( RRArbiter_0_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( RRArbiter_0_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( RRArbiter_0_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( RRArbiter_0_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  RRArbiter_2 RRArbiter_1(.clk(clk), .reset(reset),
       .io_in_1_ready( RRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( io_in_1_finish_valid ),
       .io_in_1_bits_header_src( io_in_1_finish_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_finish_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_finish_bits_payload_master_xact_id ),
       .io_in_0_ready( RRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( io_in_0_finish_valid ),
       .io_in_0_bits_header_src( io_in_0_finish_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_finish_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_finish_bits_payload_master_xact_id ),
       .io_out_ready( io_out_finish_ready ),
       .io_out_valid( RRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( RRArbiter_1_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
endmodule

module Tile(input clk, input reset,
    input  io_tilelink_acquire_ready,
    output io_tilelink_acquire_valid,
    output[1:0] io_tilelink_acquire_bits_header_src,
    output[1:0] io_tilelink_acquire_bits_header_dst,
    output[25:0] io_tilelink_acquire_bits_payload_addr,
    output[3:0] io_tilelink_acquire_bits_payload_client_xact_id,
    output[511:0] io_tilelink_acquire_bits_payload_data,
    output[2:0] io_tilelink_acquire_bits_payload_a_type,
    output[5:0] io_tilelink_acquire_bits_payload_write_mask,
    output[2:0] io_tilelink_acquire_bits_payload_subword_addr,
    output[3:0] io_tilelink_acquire_bits_payload_atomic_opcode,
    output io_tilelink_grant_ready,
    input  io_tilelink_grant_valid,
    input [1:0] io_tilelink_grant_bits_header_src,
    input [1:0] io_tilelink_grant_bits_header_dst,
    input [511:0] io_tilelink_grant_bits_payload_data,
    input [3:0] io_tilelink_grant_bits_payload_client_xact_id,
    input [3:0] io_tilelink_grant_bits_payload_master_xact_id,
    input [3:0] io_tilelink_grant_bits_payload_g_type,
    input  io_tilelink_finish_ready,
    output io_tilelink_finish_valid,
    output[1:0] io_tilelink_finish_bits_header_src,
    output[1:0] io_tilelink_finish_bits_header_dst,
    output[3:0] io_tilelink_finish_bits_payload_master_xact_id,
    output io_tilelink_probe_ready,
    input  io_tilelink_probe_valid,
    input [1:0] io_tilelink_probe_bits_header_src,
    input [1:0] io_tilelink_probe_bits_header_dst,
    input [25:0] io_tilelink_probe_bits_payload_addr,
    input [3:0] io_tilelink_probe_bits_payload_master_xact_id,
    input [1:0] io_tilelink_probe_bits_payload_p_type,
    input  io_tilelink_release_ready,
    output io_tilelink_release_valid,
    output[1:0] io_tilelink_release_bits_header_src,
    output[1:0] io_tilelink_release_bits_header_dst,
    output[25:0] io_tilelink_release_bits_payload_addr,
    output[3:0] io_tilelink_release_bits_payload_client_xact_id,
    output[3:0] io_tilelink_release_bits_payload_master_xact_id,
    output[511:0] io_tilelink_release_bits_payload_data,
    output[2:0] io_tilelink_release_bits_payload_r_type,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr
);

  wire[3:0] dcache_io_mem_finish_bits_payload_master_xact_id;
  wire[1:0] dcache_io_mem_finish_bits_header_dst;
  wire[1:0] dcache_io_mem_finish_bits_header_src;
  wire dcache_io_mem_finish_valid;
  wire dcache_io_mem_grant_ready;
  wire[3:0] dcache_io_mem_acquire_bits_payload_atomic_opcode;
  wire[2:0] dcache_io_mem_acquire_bits_payload_subword_addr;
  wire[5:0] dcache_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] dcache_io_mem_acquire_bits_payload_a_type;
  wire[511:0] dcache_io_mem_acquire_bits_payload_data;
  wire[3:0] dcache_io_mem_acquire_bits_payload_client_xact_id;
  wire[25:0] dcache_io_mem_acquire_bits_payload_addr;
  wire[1:0] dcache_io_mem_acquire_bits_header_dst;
  wire[1:0] dcache_io_mem_acquire_bits_header_src;
  wire dcache_io_mem_acquire_valid;
  wire[3:0] icache_io_mem_finish_bits_payload_master_xact_id;
  wire[1:0] icache_io_mem_finish_bits_header_dst;
  wire[1:0] icache_io_mem_finish_bits_header_src;
  wire icache_io_mem_finish_valid;
  wire icache_io_mem_grant_ready;
  wire[3:0] icache_io_mem_acquire_bits_payload_atomic_opcode;
  wire[2:0] icache_io_mem_acquire_bits_payload_subword_addr;
  wire[5:0] icache_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] icache_io_mem_acquire_bits_payload_a_type;
  wire[511:0] icache_io_mem_acquire_bits_payload_data;
  wire[3:0] icache_io_mem_acquire_bits_payload_client_xact_id;
  wire[25:0] icache_io_mem_acquire_bits_payload_addr;
  wire icache_io_mem_acquire_valid;
  wire dcache_io_cpu_ordered;
  wire[29:0] dcache_io_cpu_ptw_req_bits;
  wire dcache_io_cpu_ptw_req_valid;
  wire dcache_io_cpu_xcpt_pf_st;
  wire dcache_io_cpu_xcpt_pf_ld;
  wire dcache_io_cpu_xcpt_ma_st;
  wire dcache_io_cpu_xcpt_ma_ld;
  wire[7:0] dcache_io_cpu_replay_next_bits;
  wire dcache_io_cpu_replay_next_valid;
  wire[63:0] dcache_io_cpu_resp_bits_store_data;
  wire[43:0] dcache_io_cpu_resp_bits_addr;
  wire[3:0] dcache_io_cpu_resp_bits_cmd;
  wire[7:0] dcache_io_cpu_resp_bits_tag;
  wire[63:0] dcache_io_cpu_resp_bits_data_subword;
  wire[63:0] dcache_io_cpu_resp_bits_data;
  wire dcache_io_cpu_resp_bits_has_data;
  wire[2:0] dcache_io_cpu_resp_bits_typ;
  wire dcache_io_cpu_resp_bits_replay;
  wire dcache_io_cpu_resp_bits_nack;
  wire dcache_io_cpu_resp_valid;
  wire dcache_io_cpu_req_ready;
  wire[4:0] ptw_io_mem_req_bits_cmd;
  wire[43:0] ptw_io_mem_req_bits_addr;
  wire ptw_io_mem_req_bits_phys;
  wire[2:0] ptw_io_mem_req_bits_typ;
  wire ptw_io_mem_req_bits_kill;
  wire ptw_io_mem_req_valid;
  wire[4:0] core_io_dmem_req_bits_cmd;
  wire[7:0] core_io_dmem_req_bits_tag;
  wire[63:0] core_io_dmem_req_bits_data;
  wire[43:0] core_io_dmem_req_bits_addr;
  wire core_io_dmem_req_bits_phys;
  wire[2:0] core_io_dmem_req_bits_typ;
  wire core_io_dmem_req_bits_kill;
  wire core_io_dmem_req_valid;
  wire core_io_ptw_status_s;
  wire core_io_ptw_status_ps;
  wire core_io_ptw_status_ei;
  wire core_io_ptw_status_pei;
  wire core_io_ptw_status_ef;
  wire core_io_ptw_status_u64;
  wire core_io_ptw_status_s64;
  wire core_io_ptw_status_vm;
  wire core_io_ptw_status_er;
  wire[6:0] core_io_ptw_status_zero;
  wire[7:0] core_io_ptw_status_im;
  wire[7:0] core_io_ptw_status_ip;
  wire core_io_ptw_sret;
  wire core_io_ptw_invalidate;
  wire[31:0] core_io_ptw_ptbr;
  wire dcacheArb_io_requestor_0_ordered;
  wire dcacheArb_io_requestor_0_xcpt_pf_st;
  wire dcacheArb_io_requestor_0_xcpt_pf_ld;
  wire dcacheArb_io_requestor_0_xcpt_ma_st;
  wire dcacheArb_io_requestor_0_xcpt_ma_ld;
  wire[7:0] dcacheArb_io_requestor_0_replay_next_bits;
  wire dcacheArb_io_requestor_0_replay_next_valid;
  wire[63:0] dcacheArb_io_requestor_0_resp_bits_store_data;
  wire[43:0] dcacheArb_io_requestor_0_resp_bits_addr;
  wire[3:0] dcacheArb_io_requestor_0_resp_bits_cmd;
  wire[7:0] dcacheArb_io_requestor_0_resp_bits_tag;
  wire[63:0] dcacheArb_io_requestor_0_resp_bits_data_subword;
  wire[63:0] dcacheArb_io_requestor_0_resp_bits_data;
  wire dcacheArb_io_requestor_0_resp_bits_has_data;
  wire[2:0] dcacheArb_io_requestor_0_resp_bits_typ;
  wire dcacheArb_io_requestor_0_resp_bits_replay;
  wire dcacheArb_io_requestor_0_resp_bits_nack;
  wire dcacheArb_io_requestor_0_resp_valid;
  wire dcacheArb_io_requestor_0_req_ready;
  wire[29:0] icache_io_cpu_ptw_req_bits;
  wire icache_io_cpu_ptw_req_valid;
  wire memArb_io_in_0_finish_ready;
  wire[3:0] memArb_io_in_0_grant_bits_payload_g_type;
  wire[3:0] memArb_io_in_0_grant_bits_payload_master_xact_id;
  wire[3:0] memArb_io_in_0_grant_bits_payload_client_xact_id;
  wire[511:0] memArb_io_in_0_grant_bits_payload_data;
  wire[1:0] memArb_io_in_0_grant_bits_header_dst;
  wire[1:0] memArb_io_in_0_grant_bits_header_src;
  wire memArb_io_in_0_grant_valid;
  wire memArb_io_in_0_acquire_ready;
  wire ptw_io_requestor_1_sret;
  wire ptw_io_requestor_1_invalidate;
  wire ptw_io_requestor_1_status_s;
  wire ptw_io_requestor_1_status_ps;
  wire ptw_io_requestor_1_status_ei;
  wire ptw_io_requestor_1_status_pei;
  wire ptw_io_requestor_1_status_ef;
  wire ptw_io_requestor_1_status_u64;
  wire ptw_io_requestor_1_status_s64;
  wire ptw_io_requestor_1_status_vm;
  wire ptw_io_requestor_1_status_er;
  wire[6:0] ptw_io_requestor_1_status_zero;
  wire[7:0] ptw_io_requestor_1_status_im;
  wire[7:0] ptw_io_requestor_1_status_ip;
  wire[5:0] ptw_io_requestor_1_resp_bits_perm;
  wire[18:0] ptw_io_requestor_1_resp_bits_ppn;
  wire ptw_io_requestor_1_resp_bits_error;
  wire ptw_io_requestor_1_resp_valid;
  wire ptw_io_requestor_1_req_ready;
  wire[4:0] dcacheArb_io_mem_req_bits_cmd;
  wire[7:0] dcacheArb_io_mem_req_bits_tag;
  wire[63:0] dcacheArb_io_mem_req_bits_data;
  wire[43:0] dcacheArb_io_mem_req_bits_addr;
  wire dcacheArb_io_mem_req_bits_phys;
  wire[2:0] dcacheArb_io_mem_req_bits_typ;
  wire dcacheArb_io_mem_req_bits_kill;
  wire dcacheArb_io_mem_req_valid;
  wire memArb_io_in_1_finish_ready;
  wire[3:0] memArb_io_in_1_grant_bits_payload_g_type;
  wire[3:0] memArb_io_in_1_grant_bits_payload_master_xact_id;
  wire[3:0] memArb_io_in_1_grant_bits_payload_client_xact_id;
  wire[511:0] memArb_io_in_1_grant_bits_payload_data;
  wire[1:0] memArb_io_in_1_grant_bits_header_dst;
  wire[1:0] memArb_io_in_1_grant_bits_header_src;
  wire memArb_io_in_1_grant_valid;
  wire memArb_io_in_1_acquire_ready;
  wire core_io_imem_invalidate;
  wire ptw_io_requestor_0_sret;
  wire ptw_io_requestor_0_invalidate;
  wire ptw_io_requestor_0_status_s;
  wire ptw_io_requestor_0_status_ps;
  wire ptw_io_requestor_0_status_ei;
  wire ptw_io_requestor_0_status_pei;
  wire ptw_io_requestor_0_status_ef;
  wire ptw_io_requestor_0_status_u64;
  wire ptw_io_requestor_0_status_s64;
  wire ptw_io_requestor_0_status_vm;
  wire ptw_io_requestor_0_status_er;
  wire[6:0] ptw_io_requestor_0_status_zero;
  wire[7:0] ptw_io_requestor_0_status_im;
  wire[7:0] ptw_io_requestor_0_status_ip;
  wire[5:0] ptw_io_requestor_0_resp_bits_perm;
  wire[18:0] ptw_io_requestor_0_resp_bits_ppn;
  wire ptw_io_requestor_0_resp_bits_error;
  wire ptw_io_requestor_0_resp_valid;
  wire ptw_io_requestor_0_req_ready;
  wire core_io_imem_btb_update_bits_incorrectTarget;
  wire core_io_imem_btb_update_bits_isReturn;
  wire core_io_imem_btb_update_bits_isCall;
  wire core_io_imem_btb_update_bits_isJump;
  wire core_io_imem_btb_update_bits_taken;
  wire[42:0] core_io_imem_btb_update_bits_returnAddr;
  wire[42:0] core_io_imem_btb_update_bits_target;
  wire[42:0] core_io_imem_btb_update_bits_pc;
  wire[1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire[3:0] core_io_imem_btb_update_bits_prediction_bits_bht_index;
  wire[2:0] core_io_imem_btb_update_bits_prediction_bits_entry;
  wire[42:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire core_io_imem_btb_update_bits_prediction_bits_taken;
  wire core_io_imem_btb_update_bits_prediction_valid;
  wire core_io_imem_btb_update_valid;
  wire core_io_imem_resp_ready;
  wire[43:0] core_io_imem_req_bits_pc;
  wire core_io_imem_req_valid;
  wire dcacheArb_io_requestor_1_ordered;
  wire dcacheArb_io_requestor_1_xcpt_pf_st;
  wire dcacheArb_io_requestor_1_xcpt_pf_ld;
  wire dcacheArb_io_requestor_1_xcpt_ma_st;
  wire dcacheArb_io_requestor_1_xcpt_ma_ld;
  wire[7:0] dcacheArb_io_requestor_1_replay_next_bits;
  wire dcacheArb_io_requestor_1_replay_next_valid;
  wire[63:0] dcacheArb_io_requestor_1_resp_bits_store_data;
  wire[43:0] dcacheArb_io_requestor_1_resp_bits_addr;
  wire[3:0] dcacheArb_io_requestor_1_resp_bits_cmd;
  wire[7:0] dcacheArb_io_requestor_1_resp_bits_tag;
  wire[63:0] dcacheArb_io_requestor_1_resp_bits_data_subword;
  wire[63:0] dcacheArb_io_requestor_1_resp_bits_data;
  wire dcacheArb_io_requestor_1_resp_bits_has_data;
  wire[2:0] dcacheArb_io_requestor_1_resp_bits_typ;
  wire dcacheArb_io_requestor_1_resp_bits_replay;
  wire dcacheArb_io_requestor_1_resp_bits_nack;
  wire dcacheArb_io_requestor_1_resp_valid;
  wire dcacheArb_io_requestor_1_req_ready;
  wire[1:0] icache_io_cpu_btb_resp_bits_bht_value;
  wire[3:0] icache_io_cpu_btb_resp_bits_bht_index;
  wire[2:0] icache_io_cpu_btb_resp_bits_entry;
  wire[42:0] icache_io_cpu_btb_resp_bits_target;
  wire icache_io_cpu_btb_resp_bits_taken;
  wire icache_io_cpu_btb_resp_valid;
  wire icache_io_cpu_resp_bits_xcpt_if;
  wire icache_io_cpu_resp_bits_xcpt_ma;
  wire[31:0] icache_io_cpu_resp_bits_data;
  wire[43:0] icache_io_cpu_resp_bits_pc;
  wire icache_io_cpu_resp_valid;
  wire core_io_host_debug_stats_pcr;
  wire core_io_host_ipi_rep_ready;
  wire core_io_host_ipi_req_bits;
  wire core_io_host_ipi_req_valid;
  wire[63:0] core_io_host_pcr_rep_bits;
  wire core_io_host_pcr_rep_valid;
  wire core_io_host_pcr_req_ready;
  wire[2:0] dcache_io_mem_release_bits_payload_r_type;
  wire[511:0] dcache_io_mem_release_bits_payload_data;
  wire[3:0] dcache_io_mem_release_bits_payload_master_xact_id;
  wire[3:0] T0;
  wire[4:0] T1;
  wire[3:0] dcache_io_mem_release_bits_payload_client_xact_id;
  wire[25:0] dcache_io_mem_release_bits_payload_addr;
  wire[1:0] dcache_io_mem_release_bits_header_dst;
  wire[1:0] dcache_io_mem_release_bits_header_src;
  wire dcache_io_mem_release_valid;
  wire dcache_io_mem_probe_ready;
  wire[3:0] memArb_io_out_finish_bits_payload_master_xact_id;
  wire[1:0] memArb_io_out_finish_bits_header_dst;
  wire[1:0] memArb_io_out_finish_bits_header_src;
  wire memArb_io_out_finish_valid;
  wire memArb_io_out_grant_ready;
  wire[3:0] memArb_io_out_acquire_bits_payload_atomic_opcode;
  wire[2:0] memArb_io_out_acquire_bits_payload_subword_addr;
  wire[5:0] memArb_io_out_acquire_bits_payload_write_mask;
  wire[2:0] memArb_io_out_acquire_bits_payload_a_type;
  wire[511:0] memArb_io_out_acquire_bits_payload_data;
  wire[3:0] memArb_io_out_acquire_bits_payload_client_xact_id;
  wire[25:0] memArb_io_out_acquire_bits_payload_addr;
  wire[1:0] memArb_io_out_acquire_bits_header_dst;
  wire[1:0] memArb_io_out_acquire_bits_header_src;
  wire memArb_io_out_acquire_valid;


  assign io_host_debug_stats_pcr = core_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = core_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = core_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = core_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = core_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = core_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = core_io_host_pcr_req_ready;
  assign io_tilelink_release_bits_payload_r_type = dcache_io_mem_release_bits_payload_r_type;
  assign io_tilelink_release_bits_payload_data = dcache_io_mem_release_bits_payload_data;
  assign io_tilelink_release_bits_payload_master_xact_id = dcache_io_mem_release_bits_payload_master_xact_id;
  assign io_tilelink_release_bits_payload_client_xact_id = T0;
  assign T0 = T1[2'h3:1'h0];
  assign T1 = {dcache_io_mem_release_bits_payload_client_xact_id, 1'h0};
  assign io_tilelink_release_bits_payload_addr = dcache_io_mem_release_bits_payload_addr;
  assign io_tilelink_release_bits_header_dst = dcache_io_mem_release_bits_header_dst;
  assign io_tilelink_release_bits_header_src = dcache_io_mem_release_bits_header_src;
  assign io_tilelink_release_valid = dcache_io_mem_release_valid;
  assign io_tilelink_probe_ready = dcache_io_mem_probe_ready;
  assign io_tilelink_finish_bits_payload_master_xact_id = memArb_io_out_finish_bits_payload_master_xact_id;
  assign io_tilelink_finish_bits_header_dst = memArb_io_out_finish_bits_header_dst;
  assign io_tilelink_finish_bits_header_src = memArb_io_out_finish_bits_header_src;
  assign io_tilelink_finish_valid = memArb_io_out_finish_valid;
  assign io_tilelink_grant_ready = memArb_io_out_grant_ready;
  assign io_tilelink_acquire_bits_payload_atomic_opcode = memArb_io_out_acquire_bits_payload_atomic_opcode;
  assign io_tilelink_acquire_bits_payload_subword_addr = memArb_io_out_acquire_bits_payload_subword_addr;
  assign io_tilelink_acquire_bits_payload_write_mask = memArb_io_out_acquire_bits_payload_write_mask;
  assign io_tilelink_acquire_bits_payload_a_type = memArb_io_out_acquire_bits_payload_a_type;
  assign io_tilelink_acquire_bits_payload_data = memArb_io_out_acquire_bits_payload_data;
  assign io_tilelink_acquire_bits_payload_client_xact_id = memArb_io_out_acquire_bits_payload_client_xact_id;
  assign io_tilelink_acquire_bits_payload_addr = memArb_io_out_acquire_bits_payload_addr;
  assign io_tilelink_acquire_bits_header_dst = memArb_io_out_acquire_bits_header_dst;
  assign io_tilelink_acquire_bits_header_src = memArb_io_out_acquire_bits_header_src;
  assign io_tilelink_acquire_valid = memArb_io_out_acquire_valid;
  Core core(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( core_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( core_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( core_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( core_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( core_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( core_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( core_io_host_debug_stats_pcr ),
       .io_imem_req_valid( core_io_imem_req_valid ),
       .io_imem_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_imem_resp_ready( core_io_imem_resp_ready ),
       .io_imem_resp_valid( icache_io_cpu_resp_valid ),
       .io_imem_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_imem_resp_bits_data( icache_io_cpu_resp_bits_data ),
       .io_imem_resp_bits_xcpt_ma( icache_io_cpu_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_index( icache_io_cpu_btb_resp_bits_bht_index ),
       .io_imem_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_index( core_io_imem_btb_update_bits_prediction_bits_bht_index ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_imem_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       .io_imem_btb_update_bits_returnAddr( core_io_imem_btb_update_bits_returnAddr ),
       .io_imem_btb_update_bits_taken( core_io_imem_btb_update_bits_taken ),
       .io_imem_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isCall( core_io_imem_btb_update_bits_isCall ),
       .io_imem_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_imem_btb_update_bits_incorrectTarget( core_io_imem_btb_update_bits_incorrectTarget ),
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_imem_ptw_req_bits( icache_io_cpu_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       .io_imem_invalidate( core_io_imem_invalidate ),
       .io_dmem_req_ready( dcacheArb_io_requestor_1_req_ready ),
       .io_dmem_req_valid( core_io_dmem_req_valid ),
       .io_dmem_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_dmem_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_data( core_io_dmem_req_bits_data ),
       .io_dmem_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_dmem_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_dmem_resp_valid( dcacheArb_io_requestor_1_resp_valid ),
       .io_dmem_resp_bits_nack( dcacheArb_io_requestor_1_resp_bits_nack ),
       .io_dmem_resp_bits_replay( dcacheArb_io_requestor_1_resp_bits_replay ),
       .io_dmem_resp_bits_typ( dcacheArb_io_requestor_1_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( dcacheArb_io_requestor_1_resp_bits_has_data ),
       .io_dmem_resp_bits_data( dcacheArb_io_requestor_1_resp_bits_data ),
       .io_dmem_resp_bits_data_subword( dcacheArb_io_requestor_1_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( dcacheArb_io_requestor_1_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( dcacheArb_io_requestor_1_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( dcacheArb_io_requestor_1_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( dcacheArb_io_requestor_1_resp_bits_store_data ),
       .io_dmem_replay_next_valid( dcacheArb_io_requestor_1_replay_next_valid ),
       .io_dmem_replay_next_bits( dcacheArb_io_requestor_1_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( dcacheArb_io_requestor_1_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( dcacheArb_io_requestor_1_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( dcacheArb_io_requestor_1_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( dcacheArb_io_requestor_1_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       //.io_dmem_ptw_req_valid(  )
       //.io_dmem_ptw_req_bits(  )
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( dcacheArb_io_requestor_1_ordered ),
       .io_ptw_ptbr( core_io_ptw_ptbr ),
       .io_ptw_invalidate( core_io_ptw_invalidate ),
       .io_ptw_sret( core_io_ptw_sret ),
       .io_ptw_status_ip( core_io_ptw_status_ip ),
       .io_ptw_status_im( core_io_ptw_status_im ),
       .io_ptw_status_zero( core_io_ptw_status_zero ),
       .io_ptw_status_er( core_io_ptw_status_er ),
       .io_ptw_status_vm( core_io_ptw_status_vm ),
       .io_ptw_status_s64( core_io_ptw_status_s64 ),
       .io_ptw_status_u64( core_io_ptw_status_u64 ),
       .io_ptw_status_ef( core_io_ptw_status_ef ),
       .io_ptw_status_pei( core_io_ptw_status_pei ),
       .io_ptw_status_ei( core_io_ptw_status_ei ),
       .io_ptw_status_ps( core_io_ptw_status_ps ),
       .io_ptw_status_s( core_io_ptw_status_s )
       //.io_rocc_cmd_ready(  )
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       //.io_rocc_resp_valid(  )
       //.io_rocc_resp_bits_rd(  )
       //.io_rocc_resp_bits_data(  )
       //.io_rocc_mem_req_ready(  )
       //.io_rocc_mem_req_valid(  )
       //.io_rocc_mem_req_bits_kill(  )
       //.io_rocc_mem_req_bits_typ(  )
       //.io_rocc_mem_req_bits_phys(  )
       //.io_rocc_mem_req_bits_addr(  )
       //.io_rocc_mem_req_bits_data(  )
       //.io_rocc_mem_req_bits_tag(  )
       //.io_rocc_mem_req_bits_cmd(  )
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       //.io_rocc_mem_ptw_req_ready(  )
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       //.io_rocc_mem_ptw_resp_valid(  )
       //.io_rocc_mem_ptw_resp_bits_error(  )
       //.io_rocc_mem_ptw_resp_bits_ppn(  )
       //.io_rocc_mem_ptw_resp_bits_perm(  )
       //.io_rocc_mem_ptw_status_ip(  )
       //.io_rocc_mem_ptw_status_im(  )
       //.io_rocc_mem_ptw_status_zero(  )
       //.io_rocc_mem_ptw_status_er(  )
       //.io_rocc_mem_ptw_status_vm(  )
       //.io_rocc_mem_ptw_status_s64(  )
       //.io_rocc_mem_ptw_status_u64(  )
       //.io_rocc_mem_ptw_status_ef(  )
       //.io_rocc_mem_ptw_status_pei(  )
       //.io_rocc_mem_ptw_status_ei(  )
       //.io_rocc_mem_ptw_status_ps(  )
       //.io_rocc_mem_ptw_status_s(  )
       //.io_rocc_mem_ptw_invalidate(  )
       //.io_rocc_mem_ptw_sret(  )
       //.io_rocc_mem_ordered(  )
       //.io_rocc_busy(  )
       //.io_rocc_s(  )
       //.io_rocc_interrupt(  )
       //.io_rocc_imem_acquire_ready(  )
       //.io_rocc_imem_acquire_valid(  )
       //.io_rocc_imem_acquire_bits_header_src(  )
       //.io_rocc_imem_acquire_bits_header_dst(  )
       //.io_rocc_imem_acquire_bits_payload_addr(  )
       //.io_rocc_imem_acquire_bits_payload_client_xact_id(  )
       //.io_rocc_imem_acquire_bits_payload_data(  )
       //.io_rocc_imem_acquire_bits_payload_a_type(  )
       //.io_rocc_imem_acquire_bits_payload_write_mask(  )
       //.io_rocc_imem_acquire_bits_payload_subword_addr(  )
       //.io_rocc_imem_acquire_bits_payload_atomic_opcode(  )
       //.io_rocc_imem_grant_ready(  )
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       //.io_rocc_imem_finish_valid(  )
       //.io_rocc_imem_finish_bits_header_src(  )
       //.io_rocc_imem_finish_bits_header_dst(  )
       //.io_rocc_imem_finish_bits_payload_master_xact_id(  )
       //.io_rocc_iptw_req_ready(  )
       //.io_rocc_iptw_req_valid(  )
       //.io_rocc_iptw_req_bits(  )
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       //.io_rocc_dptw_req_valid(  )
       //.io_rocc_dptw_req_bits(  )
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       //.io_rocc_pptw_req_valid(  )
       //.io_rocc_pptw_req_bits(  )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
  );
  `ifndef SYNTHESIS
    assign core.io_dmem_ptw_req_valid = {1{$random}};
    assign core.io_dmem_ptw_req_bits = {1{$random}};
    assign core.io_rocc_cmd_ready = {1{$random}};
    assign core.io_rocc_resp_valid = {1{$random}};
    assign core.io_rocc_resp_bits_rd = {1{$random}};
    assign core.io_rocc_resp_bits_data = {2{$random}};
    assign core.io_rocc_mem_req_valid = {1{$random}};
    assign core.io_rocc_mem_req_bits_kill = {1{$random}};
    assign core.io_rocc_mem_req_bits_typ = {1{$random}};
    assign core.io_rocc_mem_req_bits_phys = {1{$random}};
    assign core.io_rocc_mem_req_bits_addr = {2{$random}};
    assign core.io_rocc_mem_req_bits_data = {2{$random}};
    assign core.io_rocc_mem_req_bits_tag = {1{$random}};
    assign core.io_rocc_mem_req_bits_cmd = {1{$random}};
    assign core.io_rocc_mem_ptw_req_ready = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_valid = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_error = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_ppn = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_perm = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ip = {1{$random}};
    assign core.io_rocc_mem_ptw_status_im = {1{$random}};
    assign core.io_rocc_mem_ptw_status_zero = {1{$random}};
    assign core.io_rocc_mem_ptw_status_er = {1{$random}};
    assign core.io_rocc_mem_ptw_status_vm = {1{$random}};
    assign core.io_rocc_mem_ptw_status_s64 = {1{$random}};
    assign core.io_rocc_mem_ptw_status_u64 = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ef = {1{$random}};
    assign core.io_rocc_mem_ptw_status_pei = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ei = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ps = {1{$random}};
    assign core.io_rocc_mem_ptw_status_s = {1{$random}};
    assign core.io_rocc_mem_ptw_invalidate = {1{$random}};
    assign core.io_rocc_mem_ptw_sret = {1{$random}};
    assign core.io_rocc_busy = {1{$random}};
    assign core.io_rocc_interrupt = {1{$random}};
    assign core.io_rocc_imem_acquire_valid = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_header_src = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_header_dst = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_addr = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_client_xact_id = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_data = {16{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_a_type = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_write_mask = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_subword_addr = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_atomic_opcode = {1{$random}};
    assign core.io_rocc_imem_grant_ready = {1{$random}};
    assign core.io_rocc_imem_finish_valid = {1{$random}};
    assign core.io_rocc_imem_finish_bits_header_src = {1{$random}};
    assign core.io_rocc_imem_finish_bits_header_dst = {1{$random}};
    assign core.io_rocc_imem_finish_bits_payload_master_xact_id = {1{$random}};
    assign core.io_rocc_iptw_req_valid = {1{$random}};
    assign core.io_rocc_iptw_req_bits = {1{$random}};
    assign core.io_rocc_dptw_req_valid = {1{$random}};
    assign core.io_rocc_dptw_req_bits = {1{$random}};
    assign core.io_rocc_pptw_req_valid = {1{$random}};
    assign core.io_rocc_pptw_req_bits = {1{$random}};
  `endif
  Frontend icache(.clk(clk), .reset(reset),
       .io_cpu_req_valid( core_io_imem_req_valid ),
       .io_cpu_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_cpu_resp_ready( core_io_imem_resp_ready ),
       .io_cpu_resp_valid( icache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_cpu_resp_bits_data( icache_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_xcpt_ma( icache_io_cpu_resp_bits_xcpt_ma ),
       .io_cpu_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_cpu_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_cpu_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_cpu_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_cpu_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_cpu_btb_resp_bits_bht_index( icache_io_cpu_btb_resp_bits_bht_index ),
       .io_cpu_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_cpu_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_cpu_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_cpu_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_cpu_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_cpu_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_cpu_btb_update_bits_prediction_bits_bht_index( core_io_imem_btb_update_bits_prediction_bits_bht_index ),
       .io_cpu_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_cpu_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_cpu_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       .io_cpu_btb_update_bits_returnAddr( core_io_imem_btb_update_bits_returnAddr ),
       .io_cpu_btb_update_bits_taken( core_io_imem_btb_update_bits_taken ),
       .io_cpu_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_cpu_btb_update_bits_isCall( core_io_imem_btb_update_bits_isCall ),
       .io_cpu_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_cpu_btb_update_bits_incorrectTarget( core_io_imem_btb_update_bits_incorrectTarget ),
       .io_cpu_ptw_req_ready( ptw_io_requestor_0_req_ready ),
       .io_cpu_ptw_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_cpu_ptw_req_bits( icache_io_cpu_ptw_req_bits ),
       .io_cpu_ptw_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_cpu_ptw_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_cpu_ptw_resp_bits_ppn( ptw_io_requestor_0_resp_bits_ppn ),
       .io_cpu_ptw_resp_bits_perm( ptw_io_requestor_0_resp_bits_perm ),
       .io_cpu_ptw_status_ip( ptw_io_requestor_0_status_ip ),
       .io_cpu_ptw_status_im( ptw_io_requestor_0_status_im ),
       .io_cpu_ptw_status_zero( ptw_io_requestor_0_status_zero ),
       .io_cpu_ptw_status_er( ptw_io_requestor_0_status_er ),
       .io_cpu_ptw_status_vm( ptw_io_requestor_0_status_vm ),
       .io_cpu_ptw_status_s64( ptw_io_requestor_0_status_s64 ),
       .io_cpu_ptw_status_u64( ptw_io_requestor_0_status_u64 ),
       .io_cpu_ptw_status_ef( ptw_io_requestor_0_status_ef ),
       .io_cpu_ptw_status_pei( ptw_io_requestor_0_status_pei ),
       .io_cpu_ptw_status_ei( ptw_io_requestor_0_status_ei ),
       .io_cpu_ptw_status_ps( ptw_io_requestor_0_status_ps ),
       .io_cpu_ptw_status_s( ptw_io_requestor_0_status_s ),
       .io_cpu_ptw_invalidate( ptw_io_requestor_0_invalidate ),
       .io_cpu_ptw_sret( ptw_io_requestor_0_sret ),
       .io_cpu_invalidate( core_io_imem_invalidate ),
       .io_mem_acquire_ready( memArb_io_in_1_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( icache_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( icache_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( icache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( memArb_io_in_1_grant_valid ),
       .io_mem_grant_bits_header_src( memArb_io_in_1_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( memArb_io_in_1_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( memArb_io_in_1_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( memArb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( memArb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( memArb_io_in_1_grant_bits_payload_g_type ),
       .io_mem_finish_ready( memArb_io_in_1_finish_ready ),
       .io_mem_finish_valid( icache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( icache_io_mem_finish_bits_payload_master_xact_id )
  );
  HellaCache dcache(.clk(clk), .reset(reset),
       .io_cpu_req_ready( dcache_io_cpu_req_ready ),
       .io_cpu_req_valid( dcacheArb_io_mem_req_valid ),
       .io_cpu_req_bits_kill( dcacheArb_io_mem_req_bits_kill ),
       .io_cpu_req_bits_typ( dcacheArb_io_mem_req_bits_typ ),
       .io_cpu_req_bits_phys( dcacheArb_io_mem_req_bits_phys ),
       .io_cpu_req_bits_addr( dcacheArb_io_mem_req_bits_addr ),
       .io_cpu_req_bits_data( dcacheArb_io_mem_req_bits_data ),
       .io_cpu_req_bits_tag( dcacheArb_io_mem_req_bits_tag ),
       .io_cpu_req_bits_cmd( dcacheArb_io_mem_req_bits_cmd ),
       .io_cpu_resp_valid( dcache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_cpu_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_cpu_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_cpu_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_cpu_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_data_subword( dcache_io_cpu_resp_bits_data_subword ),
       .io_cpu_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_cpu_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_cpu_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_cpu_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_cpu_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_cpu_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_cpu_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_cpu_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_cpu_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_cpu_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       .io_cpu_ptw_req_ready( ptw_io_requestor_1_req_ready ),
       .io_cpu_ptw_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_cpu_ptw_req_bits( dcache_io_cpu_ptw_req_bits ),
       .io_cpu_ptw_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_cpu_ptw_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_cpu_ptw_resp_bits_ppn( ptw_io_requestor_1_resp_bits_ppn ),
       .io_cpu_ptw_resp_bits_perm( ptw_io_requestor_1_resp_bits_perm ),
       .io_cpu_ptw_status_ip( ptw_io_requestor_1_status_ip ),
       .io_cpu_ptw_status_im( ptw_io_requestor_1_status_im ),
       .io_cpu_ptw_status_zero( ptw_io_requestor_1_status_zero ),
       .io_cpu_ptw_status_er( ptw_io_requestor_1_status_er ),
       .io_cpu_ptw_status_vm( ptw_io_requestor_1_status_vm ),
       .io_cpu_ptw_status_s64( ptw_io_requestor_1_status_s64 ),
       .io_cpu_ptw_status_u64( ptw_io_requestor_1_status_u64 ),
       .io_cpu_ptw_status_ef( ptw_io_requestor_1_status_ef ),
       .io_cpu_ptw_status_pei( ptw_io_requestor_1_status_pei ),
       .io_cpu_ptw_status_ei( ptw_io_requestor_1_status_ei ),
       .io_cpu_ptw_status_ps( ptw_io_requestor_1_status_ps ),
       .io_cpu_ptw_status_s( ptw_io_requestor_1_status_s ),
       .io_cpu_ptw_invalidate( ptw_io_requestor_1_invalidate ),
       .io_cpu_ptw_sret( ptw_io_requestor_1_sret ),
       .io_cpu_ordered( dcache_io_cpu_ordered ),
       .io_mem_acquire_ready( memArb_io_in_0_acquire_ready ),
       .io_mem_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_header_src( dcache_io_mem_acquire_bits_header_src ),
       .io_mem_acquire_bits_header_dst( dcache_io_mem_acquire_bits_header_dst ),
       .io_mem_acquire_bits_payload_addr( dcache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( dcache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( dcache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( dcache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( dcache_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( dcache_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( dcache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( dcache_io_mem_grant_ready ),
       .io_mem_grant_valid( memArb_io_in_0_grant_valid ),
       .io_mem_grant_bits_header_src( memArb_io_in_0_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( memArb_io_in_0_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( memArb_io_in_0_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( memArb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( memArb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( memArb_io_in_0_grant_bits_payload_g_type ),
       .io_mem_finish_ready( memArb_io_in_0_finish_ready ),
       .io_mem_finish_valid( dcache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( dcache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( dcache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( dcache_io_mem_finish_bits_payload_master_xact_id ),
       .io_mem_probe_ready( dcache_io_mem_probe_ready ),
       .io_mem_probe_valid( io_tilelink_probe_valid ),
       .io_mem_probe_bits_header_src( io_tilelink_probe_bits_header_src ),
       .io_mem_probe_bits_header_dst( io_tilelink_probe_bits_header_dst ),
       .io_mem_probe_bits_payload_addr( io_tilelink_probe_bits_payload_addr ),
       .io_mem_probe_bits_payload_master_xact_id( io_tilelink_probe_bits_payload_master_xact_id ),
       .io_mem_probe_bits_payload_p_type( io_tilelink_probe_bits_payload_p_type ),
       .io_mem_release_ready( io_tilelink_release_ready ),
       .io_mem_release_valid( dcache_io_mem_release_valid ),
       .io_mem_release_bits_header_src( dcache_io_mem_release_bits_header_src ),
       .io_mem_release_bits_header_dst( dcache_io_mem_release_bits_header_dst ),
       .io_mem_release_bits_payload_addr( dcache_io_mem_release_bits_payload_addr ),
       .io_mem_release_bits_payload_client_xact_id( dcache_io_mem_release_bits_payload_client_xact_id ),
       .io_mem_release_bits_payload_master_xact_id( dcache_io_mem_release_bits_payload_master_xact_id ),
       .io_mem_release_bits_payload_data( dcache_io_mem_release_bits_payload_data ),
       .io_mem_release_bits_payload_r_type( dcache_io_mem_release_bits_payload_r_type )
  );
  PTW ptw(.clk(clk), .reset(reset),
       .io_requestor_1_req_ready( ptw_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_requestor_1_req_bits( dcache_io_cpu_ptw_req_bits ),
       .io_requestor_1_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_requestor_1_resp_bits_ppn( ptw_io_requestor_1_resp_bits_ppn ),
       .io_requestor_1_resp_bits_perm( ptw_io_requestor_1_resp_bits_perm ),
       .io_requestor_1_status_ip( ptw_io_requestor_1_status_ip ),
       .io_requestor_1_status_im( ptw_io_requestor_1_status_im ),
       .io_requestor_1_status_zero( ptw_io_requestor_1_status_zero ),
       .io_requestor_1_status_er( ptw_io_requestor_1_status_er ),
       .io_requestor_1_status_vm( ptw_io_requestor_1_status_vm ),
       .io_requestor_1_status_s64( ptw_io_requestor_1_status_s64 ),
       .io_requestor_1_status_u64( ptw_io_requestor_1_status_u64 ),
       .io_requestor_1_status_ef( ptw_io_requestor_1_status_ef ),
       .io_requestor_1_status_pei( ptw_io_requestor_1_status_pei ),
       .io_requestor_1_status_ei( ptw_io_requestor_1_status_ei ),
       .io_requestor_1_status_ps( ptw_io_requestor_1_status_ps ),
       .io_requestor_1_status_s( ptw_io_requestor_1_status_s ),
       .io_requestor_1_invalidate( ptw_io_requestor_1_invalidate ),
       .io_requestor_1_sret( ptw_io_requestor_1_sret ),
       .io_requestor_0_req_ready( ptw_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_requestor_0_req_bits( icache_io_cpu_ptw_req_bits ),
       .io_requestor_0_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_requestor_0_resp_bits_ppn( ptw_io_requestor_0_resp_bits_ppn ),
       .io_requestor_0_resp_bits_perm( ptw_io_requestor_0_resp_bits_perm ),
       .io_requestor_0_status_ip( ptw_io_requestor_0_status_ip ),
       .io_requestor_0_status_im( ptw_io_requestor_0_status_im ),
       .io_requestor_0_status_zero( ptw_io_requestor_0_status_zero ),
       .io_requestor_0_status_er( ptw_io_requestor_0_status_er ),
       .io_requestor_0_status_vm( ptw_io_requestor_0_status_vm ),
       .io_requestor_0_status_s64( ptw_io_requestor_0_status_s64 ),
       .io_requestor_0_status_u64( ptw_io_requestor_0_status_u64 ),
       .io_requestor_0_status_ef( ptw_io_requestor_0_status_ef ),
       .io_requestor_0_status_pei( ptw_io_requestor_0_status_pei ),
       .io_requestor_0_status_ei( ptw_io_requestor_0_status_ei ),
       .io_requestor_0_status_ps( ptw_io_requestor_0_status_ps ),
       .io_requestor_0_status_s( ptw_io_requestor_0_status_s ),
       .io_requestor_0_invalidate( ptw_io_requestor_0_invalidate ),
       .io_requestor_0_sret( ptw_io_requestor_0_sret ),
       .io_mem_req_ready( dcacheArb_io_requestor_0_req_ready ),
       .io_mem_req_valid( ptw_io_mem_req_valid ),
       .io_mem_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_mem_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_mem_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_mem_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_mem_req_bits_data(  )
       //.io_mem_req_bits_tag(  )
       .io_mem_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_mem_resp_valid( dcacheArb_io_requestor_0_resp_valid ),
       .io_mem_resp_bits_nack( dcacheArb_io_requestor_0_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcacheArb_io_requestor_0_resp_bits_replay ),
       .io_mem_resp_bits_typ( dcacheArb_io_requestor_0_resp_bits_typ ),
       .io_mem_resp_bits_has_data( dcacheArb_io_requestor_0_resp_bits_has_data ),
       .io_mem_resp_bits_data( dcacheArb_io_requestor_0_resp_bits_data ),
       .io_mem_resp_bits_data_subword( dcacheArb_io_requestor_0_resp_bits_data_subword ),
       .io_mem_resp_bits_tag( dcacheArb_io_requestor_0_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcacheArb_io_requestor_0_resp_bits_cmd ),
       .io_mem_resp_bits_addr( dcacheArb_io_requestor_0_resp_bits_addr ),
       .io_mem_resp_bits_store_data( dcacheArb_io_requestor_0_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcacheArb_io_requestor_0_replay_next_valid ),
       .io_mem_replay_next_bits( dcacheArb_io_requestor_0_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcacheArb_io_requestor_0_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcacheArb_io_requestor_0_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcacheArb_io_requestor_0_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcacheArb_io_requestor_0_xcpt_pf_st ),
       //.io_mem_ptw_req_ready(  )
       //.io_mem_ptw_req_valid(  )
       //.io_mem_ptw_req_bits(  )
       //.io_mem_ptw_resp_valid(  )
       //.io_mem_ptw_resp_bits_error(  )
       //.io_mem_ptw_resp_bits_ppn(  )
       //.io_mem_ptw_resp_bits_perm(  )
       //.io_mem_ptw_status_ip(  )
       //.io_mem_ptw_status_im(  )
       //.io_mem_ptw_status_zero(  )
       //.io_mem_ptw_status_er(  )
       //.io_mem_ptw_status_vm(  )
       //.io_mem_ptw_status_s64(  )
       //.io_mem_ptw_status_u64(  )
       //.io_mem_ptw_status_ef(  )
       //.io_mem_ptw_status_pei(  )
       //.io_mem_ptw_status_ei(  )
       //.io_mem_ptw_status_ps(  )
       //.io_mem_ptw_status_s(  )
       //.io_mem_ptw_invalidate(  )
       //.io_mem_ptw_sret(  )
       .io_mem_ordered( dcacheArb_io_requestor_0_ordered ),
       .io_dpath_ptbr( core_io_ptw_ptbr ),
       .io_dpath_invalidate( core_io_ptw_invalidate ),
       .io_dpath_sret( core_io_ptw_sret ),
       .io_dpath_status_ip( core_io_ptw_status_ip ),
       .io_dpath_status_im( core_io_ptw_status_im ),
       .io_dpath_status_zero( core_io_ptw_status_zero ),
       .io_dpath_status_er( core_io_ptw_status_er ),
       .io_dpath_status_vm( core_io_ptw_status_vm ),
       .io_dpath_status_s64( core_io_ptw_status_s64 ),
       .io_dpath_status_u64( core_io_ptw_status_u64 ),
       .io_dpath_status_ef( core_io_ptw_status_ef ),
       .io_dpath_status_pei( core_io_ptw_status_pei ),
       .io_dpath_status_ei( core_io_ptw_status_ei ),
       .io_dpath_status_ps( core_io_ptw_status_ps ),
       .io_dpath_status_s( core_io_ptw_status_s )
  );
  HellaCacheArbiter dcacheArb(.clk(clk),
       .io_requestor_1_req_ready( dcacheArb_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( core_io_dmem_req_valid ),
       .io_requestor_1_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_requestor_1_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_requestor_1_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_requestor_1_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_requestor_1_req_bits_data( core_io_dmem_req_bits_data ),
       .io_requestor_1_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_requestor_1_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_requestor_1_resp_valid( dcacheArb_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_nack( dcacheArb_io_requestor_1_resp_bits_nack ),
       .io_requestor_1_resp_bits_replay( dcacheArb_io_requestor_1_resp_bits_replay ),
       .io_requestor_1_resp_bits_typ( dcacheArb_io_requestor_1_resp_bits_typ ),
       .io_requestor_1_resp_bits_has_data( dcacheArb_io_requestor_1_resp_bits_has_data ),
       .io_requestor_1_resp_bits_data( dcacheArb_io_requestor_1_resp_bits_data ),
       .io_requestor_1_resp_bits_data_subword( dcacheArb_io_requestor_1_resp_bits_data_subword ),
       .io_requestor_1_resp_bits_tag( dcacheArb_io_requestor_1_resp_bits_tag ),
       .io_requestor_1_resp_bits_cmd( dcacheArb_io_requestor_1_resp_bits_cmd ),
       .io_requestor_1_resp_bits_addr( dcacheArb_io_requestor_1_resp_bits_addr ),
       .io_requestor_1_resp_bits_store_data( dcacheArb_io_requestor_1_resp_bits_store_data ),
       .io_requestor_1_replay_next_valid( dcacheArb_io_requestor_1_replay_next_valid ),
       .io_requestor_1_replay_next_bits( dcacheArb_io_requestor_1_replay_next_bits ),
       .io_requestor_1_xcpt_ma_ld( dcacheArb_io_requestor_1_xcpt_ma_ld ),
       .io_requestor_1_xcpt_ma_st( dcacheArb_io_requestor_1_xcpt_ma_st ),
       .io_requestor_1_xcpt_pf_ld( dcacheArb_io_requestor_1_xcpt_pf_ld ),
       .io_requestor_1_xcpt_pf_st( dcacheArb_io_requestor_1_xcpt_pf_st ),
       //.io_requestor_1_ptw_req_ready(  )
       //.io_requestor_1_ptw_req_valid(  )
       //.io_requestor_1_ptw_req_bits(  )
       //.io_requestor_1_ptw_resp_valid(  )
       //.io_requestor_1_ptw_resp_bits_error(  )
       //.io_requestor_1_ptw_resp_bits_ppn(  )
       //.io_requestor_1_ptw_resp_bits_perm(  )
       //.io_requestor_1_ptw_status_ip(  )
       //.io_requestor_1_ptw_status_im(  )
       //.io_requestor_1_ptw_status_zero(  )
       //.io_requestor_1_ptw_status_er(  )
       //.io_requestor_1_ptw_status_vm(  )
       //.io_requestor_1_ptw_status_s64(  )
       //.io_requestor_1_ptw_status_u64(  )
       //.io_requestor_1_ptw_status_ef(  )
       //.io_requestor_1_ptw_status_pei(  )
       //.io_requestor_1_ptw_status_ei(  )
       //.io_requestor_1_ptw_status_ps(  )
       //.io_requestor_1_ptw_status_s(  )
       //.io_requestor_1_ptw_invalidate(  )
       //.io_requestor_1_ptw_sret(  )
       .io_requestor_1_ordered( dcacheArb_io_requestor_1_ordered ),
       .io_requestor_0_req_ready( dcacheArb_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( ptw_io_mem_req_valid ),
       .io_requestor_0_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_requestor_0_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_requestor_0_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_requestor_0_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_requestor_0_req_bits_data(  )
       //.io_requestor_0_req_bits_tag(  )
       .io_requestor_0_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_requestor_0_resp_valid( dcacheArb_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_nack( dcacheArb_io_requestor_0_resp_bits_nack ),
       .io_requestor_0_resp_bits_replay( dcacheArb_io_requestor_0_resp_bits_replay ),
       .io_requestor_0_resp_bits_typ( dcacheArb_io_requestor_0_resp_bits_typ ),
       .io_requestor_0_resp_bits_has_data( dcacheArb_io_requestor_0_resp_bits_has_data ),
       .io_requestor_0_resp_bits_data( dcacheArb_io_requestor_0_resp_bits_data ),
       .io_requestor_0_resp_bits_data_subword( dcacheArb_io_requestor_0_resp_bits_data_subword ),
       .io_requestor_0_resp_bits_tag( dcacheArb_io_requestor_0_resp_bits_tag ),
       .io_requestor_0_resp_bits_cmd( dcacheArb_io_requestor_0_resp_bits_cmd ),
       .io_requestor_0_resp_bits_addr( dcacheArb_io_requestor_0_resp_bits_addr ),
       .io_requestor_0_resp_bits_store_data( dcacheArb_io_requestor_0_resp_bits_store_data ),
       .io_requestor_0_replay_next_valid( dcacheArb_io_requestor_0_replay_next_valid ),
       .io_requestor_0_replay_next_bits( dcacheArb_io_requestor_0_replay_next_bits ),
       .io_requestor_0_xcpt_ma_ld( dcacheArb_io_requestor_0_xcpt_ma_ld ),
       .io_requestor_0_xcpt_ma_st( dcacheArb_io_requestor_0_xcpt_ma_st ),
       .io_requestor_0_xcpt_pf_ld( dcacheArb_io_requestor_0_xcpt_pf_ld ),
       .io_requestor_0_xcpt_pf_st( dcacheArb_io_requestor_0_xcpt_pf_st ),
       //.io_requestor_0_ptw_req_ready(  )
       //.io_requestor_0_ptw_req_valid(  )
       //.io_requestor_0_ptw_req_bits(  )
       //.io_requestor_0_ptw_resp_valid(  )
       //.io_requestor_0_ptw_resp_bits_error(  )
       //.io_requestor_0_ptw_resp_bits_ppn(  )
       //.io_requestor_0_ptw_resp_bits_perm(  )
       //.io_requestor_0_ptw_status_ip(  )
       //.io_requestor_0_ptw_status_im(  )
       //.io_requestor_0_ptw_status_zero(  )
       //.io_requestor_0_ptw_status_er(  )
       //.io_requestor_0_ptw_status_vm(  )
       //.io_requestor_0_ptw_status_s64(  )
       //.io_requestor_0_ptw_status_u64(  )
       //.io_requestor_0_ptw_status_ef(  )
       //.io_requestor_0_ptw_status_pei(  )
       //.io_requestor_0_ptw_status_ei(  )
       //.io_requestor_0_ptw_status_ps(  )
       //.io_requestor_0_ptw_status_s(  )
       //.io_requestor_0_ptw_invalidate(  )
       //.io_requestor_0_ptw_sret(  )
       .io_requestor_0_ordered( dcacheArb_io_requestor_0_ordered ),
       .io_mem_req_ready( dcache_io_cpu_req_ready ),
       .io_mem_req_valid( dcacheArb_io_mem_req_valid ),
       .io_mem_req_bits_kill( dcacheArb_io_mem_req_bits_kill ),
       .io_mem_req_bits_typ( dcacheArb_io_mem_req_bits_typ ),
       .io_mem_req_bits_phys( dcacheArb_io_mem_req_bits_phys ),
       .io_mem_req_bits_addr( dcacheArb_io_mem_req_bits_addr ),
       .io_mem_req_bits_data( dcacheArb_io_mem_req_bits_data ),
       .io_mem_req_bits_tag( dcacheArb_io_mem_req_bits_tag ),
       .io_mem_req_bits_cmd( dcacheArb_io_mem_req_bits_cmd ),
       .io_mem_resp_valid( dcache_io_cpu_resp_valid ),
       .io_mem_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_mem_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_mem_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_mem_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_mem_resp_bits_data_subword( dcache_io_cpu_resp_bits_data_subword ),
       .io_mem_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_mem_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_mem_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_mem_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       //.io_mem_ptw_req_ready(  )
       .io_mem_ptw_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_mem_ptw_req_bits( dcache_io_cpu_ptw_req_bits ),
       //.io_mem_ptw_resp_valid(  )
       //.io_mem_ptw_resp_bits_error(  )
       //.io_mem_ptw_resp_bits_ppn(  )
       //.io_mem_ptw_resp_bits_perm(  )
       //.io_mem_ptw_status_ip(  )
       //.io_mem_ptw_status_im(  )
       //.io_mem_ptw_status_zero(  )
       //.io_mem_ptw_status_er(  )
       //.io_mem_ptw_status_vm(  )
       //.io_mem_ptw_status_s64(  )
       //.io_mem_ptw_status_u64(  )
       //.io_mem_ptw_status_ef(  )
       //.io_mem_ptw_status_pei(  )
       //.io_mem_ptw_status_ei(  )
       //.io_mem_ptw_status_ps(  )
       //.io_mem_ptw_status_s(  )
       //.io_mem_ptw_invalidate(  )
       //.io_mem_ptw_sret(  )
       .io_mem_ordered( dcache_io_cpu_ordered )
  );
  `ifndef SYNTHESIS
    assign dcacheArb.io_requestor_0_req_bits_data = {2{$random}};
    assign dcacheArb.io_requestor_0_req_bits_tag = {1{$random}};
  `endif
  UncachedTileLinkIOArbiterThatAppendsArbiterId memArb(.clk(clk), .reset(reset),
       .io_in_1_acquire_ready( memArb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_in_1_acquire_bits_header_src(  )
       //.io_in_1_acquire_bits_header_dst(  )
       .io_in_1_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_in_1_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_in_1_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_in_1_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_in_1_acquire_bits_payload_write_mask( icache_io_mem_acquire_bits_payload_write_mask ),
       .io_in_1_acquire_bits_payload_subword_addr( icache_io_mem_acquire_bits_payload_subword_addr ),
       .io_in_1_acquire_bits_payload_atomic_opcode( icache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_in_1_grant_ready( icache_io_mem_grant_ready ),
       .io_in_1_grant_valid( memArb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_header_src( memArb_io_in_1_grant_bits_header_src ),
       .io_in_1_grant_bits_header_dst( memArb_io_in_1_grant_bits_header_dst ),
       .io_in_1_grant_bits_payload_data( memArb_io_in_1_grant_bits_payload_data ),
       .io_in_1_grant_bits_payload_client_xact_id( memArb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_in_1_grant_bits_payload_master_xact_id( memArb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_in_1_grant_bits_payload_g_type( memArb_io_in_1_grant_bits_payload_g_type ),
       .io_in_1_finish_ready( memArb_io_in_1_finish_ready ),
       .io_in_1_finish_valid( icache_io_mem_finish_valid ),
       .io_in_1_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_in_1_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_in_1_finish_bits_payload_master_xact_id( icache_io_mem_finish_bits_payload_master_xact_id ),
       .io_in_0_acquire_ready( memArb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_in_0_acquire_bits_header_src( dcache_io_mem_acquire_bits_header_src ),
       .io_in_0_acquire_bits_header_dst( dcache_io_mem_acquire_bits_header_dst ),
       .io_in_0_acquire_bits_payload_addr( dcache_io_mem_acquire_bits_payload_addr ),
       .io_in_0_acquire_bits_payload_client_xact_id( dcache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_in_0_acquire_bits_payload_data( dcache_io_mem_acquire_bits_payload_data ),
       .io_in_0_acquire_bits_payload_a_type( dcache_io_mem_acquire_bits_payload_a_type ),
       .io_in_0_acquire_bits_payload_write_mask( dcache_io_mem_acquire_bits_payload_write_mask ),
       .io_in_0_acquire_bits_payload_subword_addr( dcache_io_mem_acquire_bits_payload_subword_addr ),
       .io_in_0_acquire_bits_payload_atomic_opcode( dcache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_in_0_grant_ready( dcache_io_mem_grant_ready ),
       .io_in_0_grant_valid( memArb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_header_src( memArb_io_in_0_grant_bits_header_src ),
       .io_in_0_grant_bits_header_dst( memArb_io_in_0_grant_bits_header_dst ),
       .io_in_0_grant_bits_payload_data( memArb_io_in_0_grant_bits_payload_data ),
       .io_in_0_grant_bits_payload_client_xact_id( memArb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_in_0_grant_bits_payload_master_xact_id( memArb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_in_0_grant_bits_payload_g_type( memArb_io_in_0_grant_bits_payload_g_type ),
       .io_in_0_finish_ready( memArb_io_in_0_finish_ready ),
       .io_in_0_finish_valid( dcache_io_mem_finish_valid ),
       .io_in_0_finish_bits_header_src( dcache_io_mem_finish_bits_header_src ),
       .io_in_0_finish_bits_header_dst( dcache_io_mem_finish_bits_header_dst ),
       .io_in_0_finish_bits_payload_master_xact_id( dcache_io_mem_finish_bits_payload_master_xact_id ),
       .io_out_acquire_ready( io_tilelink_acquire_ready ),
       .io_out_acquire_valid( memArb_io_out_acquire_valid ),
       .io_out_acquire_bits_header_src( memArb_io_out_acquire_bits_header_src ),
       .io_out_acquire_bits_header_dst( memArb_io_out_acquire_bits_header_dst ),
       .io_out_acquire_bits_payload_addr( memArb_io_out_acquire_bits_payload_addr ),
       .io_out_acquire_bits_payload_client_xact_id( memArb_io_out_acquire_bits_payload_client_xact_id ),
       .io_out_acquire_bits_payload_data( memArb_io_out_acquire_bits_payload_data ),
       .io_out_acquire_bits_payload_a_type( memArb_io_out_acquire_bits_payload_a_type ),
       .io_out_acquire_bits_payload_write_mask( memArb_io_out_acquire_bits_payload_write_mask ),
       .io_out_acquire_bits_payload_subword_addr( memArb_io_out_acquire_bits_payload_subword_addr ),
       .io_out_acquire_bits_payload_atomic_opcode( memArb_io_out_acquire_bits_payload_atomic_opcode ),
       .io_out_grant_ready( memArb_io_out_grant_ready ),
       .io_out_grant_valid( io_tilelink_grant_valid ),
       .io_out_grant_bits_header_src( io_tilelink_grant_bits_header_src ),
       .io_out_grant_bits_header_dst( io_tilelink_grant_bits_header_dst ),
       .io_out_grant_bits_payload_data( io_tilelink_grant_bits_payload_data ),
       .io_out_grant_bits_payload_client_xact_id( io_tilelink_grant_bits_payload_client_xact_id ),
       .io_out_grant_bits_payload_master_xact_id( io_tilelink_grant_bits_payload_master_xact_id ),
       .io_out_grant_bits_payload_g_type( io_tilelink_grant_bits_payload_g_type ),
       .io_out_finish_ready( io_tilelink_finish_ready ),
       .io_out_finish_valid( memArb_io_out_finish_valid ),
       .io_out_finish_bits_header_src( memArb_io_out_finish_bits_header_src ),
       .io_out_finish_bits_header_dst( memArb_io_out_finish_bits_header_dst ),
       .io_out_finish_bits_payload_master_xact_id( memArb_io_out_finish_bits_payload_master_xact_id )
  );
  `ifndef SYNTHESIS
    assign memArb.io_in_1_acquire_bits_header_src = {1{$random}};
    assign memArb.io_in_1_acquire_bits_header_dst = {1{$random}};
  `endif
endmodule

module Queue_2(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [3:0] io_enq_bits_client_xact_id,
    input [511:0] io_enq_bits_data,
    input [2:0] io_enq_bits_a_type,
    input [5:0] io_enq_bits_write_mask,
    input [2:0] io_enq_bits_subword_addr,
    input [3:0] io_enq_bits_atomic_opcode,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[3:0] io_deq_bits_client_xact_id,
    output[511:0] io_deq_bits_data,
    output[2:0] io_deq_bits_a_type,
    output[5:0] io_deq_bits_write_mask,
    output[2:0] io_deq_bits_subword_addr,
    output[3:0] io_deq_bits_atomic_opcode,
    output io_count
);

  wire T0;
  wire[1:0] T1;
  reg  maybe_full;
  wire T2;
  wire T3;
  wire do_enq;
  wire T4;
  wire do_flow;
  wire T5;
  wire T6;
  wire do_deq;
  wire T7;
  wire T8;
  wire[3:0] T9;
  wire[557:0] T10;
  wire[15:0] T11;
  wire[6:0] T12;
  wire[3:0] T13;
  wire[557:0] T14;
  reg [557:0] ram [0:0];
  wire[557:0] T15;
  wire[557:0] T16;
  wire[557:0] T17;
  wire[15:0] T18;
  wire[6:0] T19;
  wire[8:0] T20;
  wire[541:0] T21;
  wire[515:0] T22;
  wire[2:0] T23;
  wire[8:0] T24;
  wire[5:0] T25;
  wire[2:0] T26;
  wire[541:0] T27;
  wire[515:0] T28;
  wire[511:0] T29;
  wire[3:0] T30;
  wire[25:0] T31;
  wire[2:0] T32;
  wire[5:0] T33;
  wire[2:0] T34;
  wire[511:0] T35;
  wire[3:0] T36;
  wire[25:0] T37;
  wire T38;
  wire empty;
  wire T39;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {18{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = T1[1'h0:1'h0];
  assign T1 = {maybe_full, 1'h0};
  assign T2 = reset ? 1'h0 : T3;
  assign T3 = T6 ? do_enq : maybe_full;
  assign do_enq = T5 & T4;
  assign T4 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T5 = io_enq_ready & io_enq_valid;
  assign T6 = do_enq != do_deq;
  assign do_deq = T8 & T7;
  assign T7 = do_flow ^ 1'h1;
  assign T8 = io_deq_ready & io_deq_valid;
  assign io_deq_bits_atomic_opcode = T9;
  assign T9 = T10[2'h3:1'h0];
  assign T10 = {T27, T11};
  assign T11 = {T24, T12};
  assign T12 = {T23, T13};
  assign T13 = T14[2'h3:1'h0];
  assign T14 = ram[1'h0];
  always @(posedge clk)
    if (do_enq)
      ram[1'h0] <= T16;
  assign T16 = T17;
  assign T17 = {T21, T18};
  assign T18 = {T20, T19};
  assign T19 = {io_enq_bits_subword_addr, io_enq_bits_atomic_opcode};
  assign T20 = {io_enq_bits_a_type, io_enq_bits_write_mask};
  assign T21 = {io_enq_bits_addr, T22};
  assign T22 = {io_enq_bits_client_xact_id, io_enq_bits_data};
  assign T23 = T14[3'h6:3'h4];
  assign T24 = {T26, T25};
  assign T25 = T14[4'hc:3'h7];
  assign T26 = T14[4'hf:4'hd];
  assign T27 = {T31, T28};
  assign T28 = {T30, T29};
  assign T29 = T14[10'h20f:5'h10];
  assign T30 = T14[10'h213:10'h210];
  assign T31 = T14[10'h22d:10'h214];
  assign io_deq_bits_subword_addr = T32;
  assign T32 = T10[3'h6:3'h4];
  assign io_deq_bits_write_mask = T33;
  assign T33 = T10[4'hc:3'h7];
  assign io_deq_bits_a_type = T34;
  assign T34 = T10[4'hf:4'hd];
  assign io_deq_bits_data = T35;
  assign T35 = T10[10'h20f:5'h10];
  assign io_deq_bits_client_xact_id = T36;
  assign T36 = T10[10'h213:10'h210];
  assign io_deq_bits_addr = T37;
  assign T37 = T10[10'h22d:10'h214];
  assign io_deq_valid = T38;
  assign T38 = empty ^ 1'h1;
  assign empty = maybe_full ^ 1'h1;
  assign io_enq_ready = T39;
  assign T39 = maybe_full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T6) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module HTIF(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    output io_cpu_0_reset,
    //output io_cpu_0_id
    input  io_cpu_0_pcr_req_ready,
    output io_cpu_0_pcr_req_valid,
    output io_cpu_0_pcr_req_bits_rw,
    output[4:0] io_cpu_0_pcr_req_bits_addr,
    output[63:0] io_cpu_0_pcr_req_bits_data,
    output io_cpu_0_pcr_rep_ready,
    input  io_cpu_0_pcr_rep_valid,
    input [63:0] io_cpu_0_pcr_rep_bits,
    output io_cpu_0_ipi_req_ready,
    input  io_cpu_0_ipi_req_valid,
    input  io_cpu_0_ipi_req_bits,
    input  io_cpu_0_ipi_rep_ready,
    output io_cpu_0_ipi_rep_valid,
    //output io_cpu_0_ipi_rep_bits
    input  io_cpu_0_debug_stats_pcr,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[1:0] io_mem_acquire_bits_header_src,
    output[1:0] io_mem_acquire_bits_header_dst,
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[3:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [3:0] io_mem_grant_bits_payload_client_xact_id,
    input [3:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    //output[1:0] io_mem_finish_bits_header_src
    output[1:0] io_mem_finish_bits_header_dst,
    output[3:0] io_mem_finish_bits_payload_master_xact_id,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [1:0] io_mem_probe_bits_header_src,
    input [1:0] io_mem_probe_bits_header_dst,
    input [25:0] io_mem_probe_bits_payload_addr,
    input [3:0] io_mem_probe_bits_payload_master_xact_id,
    input [1:0] io_mem_probe_bits_payload_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    //output[1:0] io_mem_release_bits_header_src
    //output[1:0] io_mem_release_bits_header_dst
    output[25:0] io_mem_release_bits_payload_addr,
    output[3:0] io_mem_release_bits_payload_client_xact_id,
    output[3:0] io_mem_release_bits_payload_master_xact_id,
    output[511:0] io_mem_release_bits_payload_data,
    output[2:0] io_mem_release_bits_payload_r_type,
    input [63:0] io_scr_rdata_63,
    input [63:0] io_scr_rdata_62,
    input [63:0] io_scr_rdata_61,
    input [63:0] io_scr_rdata_60,
    input [63:0] io_scr_rdata_59,
    input [63:0] io_scr_rdata_58,
    input [63:0] io_scr_rdata_57,
    input [63:0] io_scr_rdata_56,
    input [63:0] io_scr_rdata_55,
    input [63:0] io_scr_rdata_54,
    input [63:0] io_scr_rdata_53,
    input [63:0] io_scr_rdata_52,
    input [63:0] io_scr_rdata_51,
    input [63:0] io_scr_rdata_50,
    input [63:0] io_scr_rdata_49,
    input [63:0] io_scr_rdata_48,
    input [63:0] io_scr_rdata_47,
    input [63:0] io_scr_rdata_46,
    input [63:0] io_scr_rdata_45,
    input [63:0] io_scr_rdata_44,
    input [63:0] io_scr_rdata_43,
    input [63:0] io_scr_rdata_42,
    input [63:0] io_scr_rdata_41,
    input [63:0] io_scr_rdata_40,
    input [63:0] io_scr_rdata_39,
    input [63:0] io_scr_rdata_38,
    input [63:0] io_scr_rdata_37,
    input [63:0] io_scr_rdata_36,
    input [63:0] io_scr_rdata_35,
    input [63:0] io_scr_rdata_34,
    input [63:0] io_scr_rdata_33,
    input [63:0] io_scr_rdata_32,
    input [63:0] io_scr_rdata_31,
    input [63:0] io_scr_rdata_30,
    input [63:0] io_scr_rdata_29,
    input [63:0] io_scr_rdata_28,
    input [63:0] io_scr_rdata_27,
    input [63:0] io_scr_rdata_26,
    input [63:0] io_scr_rdata_25,
    input [63:0] io_scr_rdata_24,
    input [63:0] io_scr_rdata_23,
    input [63:0] io_scr_rdata_22,
    input [63:0] io_scr_rdata_21,
    input [63:0] io_scr_rdata_20,
    input [63:0] io_scr_rdata_19,
    input [63:0] io_scr_rdata_18,
    input [63:0] io_scr_rdata_17,
    input [63:0] io_scr_rdata_16,
    input [63:0] io_scr_rdata_15,
    input [63:0] io_scr_rdata_14,
    input [63:0] io_scr_rdata_13,
    input [63:0] io_scr_rdata_12,
    input [63:0] io_scr_rdata_11,
    input [63:0] io_scr_rdata_10,
    input [63:0] io_scr_rdata_9,
    input [63:0] io_scr_rdata_8,
    input [63:0] io_scr_rdata_7,
    input [63:0] io_scr_rdata_6,
    input [63:0] io_scr_rdata_5,
    input [63:0] io_scr_rdata_4,
    input [63:0] io_scr_rdata_3,
    input [63:0] io_scr_rdata_2,
    //input [63:0] io_scr_rdata_1
    //input [63:0] io_scr_rdata_0
    output io_scr_wen,
    output[5:0] io_scr_waddr,
    output[63:0] io_scr_wdata
);

  wire[3:0] T0;
  wire[557:0] T1;
  wire[557:0] T2;
  wire[15:0] T3;
  wire[6:0] T4;
  wire[3:0] T5;
  wire[2:0] T6;
  wire[8:0] T7;
  wire[5:0] T8;
  wire[2:0] T9;
  wire[541:0] T10;
  wire[515:0] T11;
  wire[511:0] T12;
  wire[3:0] T13;
  wire[25:0] T14;
  wire[25:0] T15;
  wire[36:0] init_addr;
  wire[39:0] T16;
  reg [39:0] addr;
  wire[39:0] T17;
  wire[39:0] T18;
  wire[39:0] T19;
  wire[63:0] rx_shifter_in;
  wire[47:0] T20;
  reg [63:0] rx_shifter;
  wire[63:0] T21;
  wire T22;
  wire T23;
  wire T24;
  reg [14:0] rx_count;
  wire[14:0] T25;
  wire[14:0] T26;
  wire[14:0] T27;
  wire[14:0] T28;
  wire T29;
  wire T30;
  wire[12:0] T31;
  wire[11:0] tx_size;
  reg [11:0] size;
  wire[11:0] T32;
  wire[11:0] T33;
  wire T34;
  wire T35;
  wire T36;
  reg [3:0] cmd;
  wire[3:0] T37;
  wire[3:0] T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire nack;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire bad_mem_packet;
  wire T48;
  wire[2:0] T49;
  wire T50;
  wire[2:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire[12:0] T55;
  reg [14:0] tx_count;
  wire[14:0] T56;
  wire[14:0] T57;
  wire[14:0] T58;
  wire[14:0] T59;
  wire T60;
  wire T61;
  wire tx_done;
  wire T62;
  wire T63;
  wire T64;
  wire[2:0] packet_ram_raddr;
  wire[2:0] T65;
  wire T66;
  wire T67;
  wire[12:0] T68;
  wire T69;
  wire T70;
  wire[1:0] T71;
  wire T72;
  reg [3:0] state;
  wire[3:0] T73;
  wire[3:0] T74;
  wire[3:0] T75;
  wire[3:0] T76;
  wire[3:0] T77;
  wire[3:0] T78;
  wire[3:0] T79;
  wire[3:0] T80;
  wire[3:0] T81;
  wire[3:0] T82;
  wire[3:0] T83;
  wire[3:0] T84;
  wire[3:0] T85;
  wire[3:0] T86;
  wire[3:0] T87;
  wire T88;
  wire T89;
  wire[3:0] rx_cmd;
  wire T90;
  wire[12:0] rx_word_count;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire rx_done;
  wire T95;
  wire T96;
  wire T97;
  wire[2:0] T98;
  wire T99;
  wire[12:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire rx_word_done;
  wire T105;
  wire[1:0] T106;
  wire T107;
  wire T108;
  wire acq_q_io_enq_ready;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  reg  mem_acked;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire[3:0] T120;
  wire T121;
  wire T122;
  reg [8:0] pos;
  wire[8:0] T123;
  wire[8:0] T124;
  wire[8:0] T125;
  wire[8:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire[3:0] T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire[4:0] T137;
  wire T138;
  wire T139;
  wire[1:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[39:0] T145;
  wire[557:0] T146;
  wire[15:0] T147;
  wire[6:0] T148;
  wire[3:0] T149;
  wire[2:0] T150;
  wire[8:0] T151;
  wire[5:0] T152;
  wire[2:0] T153;
  wire[541:0] T154;
  wire[515:0] T155;
  wire[511:0] T156;
  wire[3:0] T157;
  wire[25:0] T158;
  wire[25:0] T159;
  wire T160;
  wire[2:0] T161;
  wire[5:0] T162;
  wire[2:0] T163;
  wire[511:0] T164;
  wire[3:0] T165;
  wire[25:0] T166;
  wire T167;
  wire T168;
  wire T169;
  wire[63:0] T170;
  reg [63:0] packet_ram_0 [7:0], packet_ram_1 [7:0], packet_ram_2 [7:0], packet_ram_3 [7:0], packet_ram_4 [7:0], packet_ram_5 [7:0], packet_ram_6 [7:0], packet_ram_7 [7:0], packet_ram_8 [7:0];
  wire[63:0] T171;
  wire[63:0] T172;
  wire T173;
  wire T174;
  wire[63:0] T175;
  wire[63:0] T176;
  wire T177;
  wire T178;
  wire[63:0] T179;
  wire[63:0] T180;
  wire T181;
  wire T182;
  wire[63:0] T183;
  wire[63:0] T184;
  wire T185;
  wire T186;
  wire[63:0] T187;
  wire[63:0] T188;
  wire T189;
  wire T190;
  wire[63:0] T191;
  wire[63:0] T192;
  wire T193;
  wire T194;
  wire[63:0] T195;
  wire[63:0] T196;
  wire T197;
  wire T198;
  wire[63:0] T199;
  wire[63:0] T200;
  wire T201;
  wire T202;
  wire[63:0] T203;
  wire T204;
  wire[2:0] T205;
  wire[2:0] T206;
  wire[5:0] T207;
  wire[5:0] T208;
  wire T209;
  wire T210;
  reg [3:0] mem_gxid;
  wire[3:0] T211;
  reg [1:0] mem_gsrc;
  wire[1:0] T212;
  wire T213;
  reg  mem_needs_ack;
  wire T214;
  wire T215;
  wire T216;
  wire[3:0] acq_q_io_deq_bits_atomic_opcode;
  wire[2:0] acq_q_io_deq_bits_subword_addr;
  wire[5:0] acq_q_io_deq_bits_write_mask;
  wire[2:0] acq_q_io_deq_bits_a_type;
  wire[511:0] mem_req_data;
  wire[447:0] T217;
  wire[383:0] T218;
  wire[319:0] T219;
  wire[255:0] T220;
  wire[191:0] T221;
  wire[127:0] T222;
  wire[63:0] T223;
  wire[63:0] T224;
  wire[63:0] T225;
  wire[63:0] T226;
  wire[63:0] T227;
  wire[63:0] T228;
  wire[63:0] T229;
  wire[63:0] T230;
  wire[3:0] acq_q_io_deq_bits_client_xact_id;
  wire[25:0] acq_q_io_deq_bits_addr;
  wire acq_q_io_deq_valid;
  reg  R231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  reg  R242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[15:0] T248;
  wire[63:0] T249;
  wire[5:0] T250;
  wire[1:0] T251;
  wire[63:0] tx_data;
  wire[63:0] T252;
  wire[63:0] T253;
  reg [63:0] pcrReadData;
  wire[63:0] T254;
  wire[63:0] T255;
  wire[63:0] T256;
  wire[63:0] T257;
  wire[63:0] T258;
  wire[63:0] T259;
  wire[63:0] T260;
  wire[63:0] T261;
  wire[63:0] T262;
  wire[63:0] T263;
  wire[63:0] scr_rdata_0;
  wire[63:0] scr_rdata_1;
  wire T264;
  wire[5:0] T265;
  wire[63:0] T266;
  wire[63:0] scr_rdata_2;
  wire[63:0] scr_rdata_3;
  wire T267;
  wire T268;
  wire[63:0] T269;
  wire[63:0] T270;
  wire[63:0] scr_rdata_4;
  wire[63:0] scr_rdata_5;
  wire T271;
  wire[63:0] T272;
  wire[63:0] scr_rdata_6;
  wire[63:0] scr_rdata_7;
  wire T273;
  wire T274;
  wire T275;
  wire[63:0] T276;
  wire[63:0] T277;
  wire[63:0] T278;
  wire[63:0] scr_rdata_8;
  wire[63:0] scr_rdata_9;
  wire T279;
  wire[63:0] T280;
  wire[63:0] scr_rdata_10;
  wire[63:0] scr_rdata_11;
  wire T281;
  wire T282;
  wire[63:0] T283;
  wire[63:0] T284;
  wire[63:0] scr_rdata_12;
  wire[63:0] scr_rdata_13;
  wire T285;
  wire[63:0] T286;
  wire[63:0] scr_rdata_14;
  wire[63:0] scr_rdata_15;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire[63:0] T291;
  wire[63:0] T292;
  wire[63:0] T293;
  wire[63:0] T294;
  wire[63:0] scr_rdata_16;
  wire[63:0] scr_rdata_17;
  wire T295;
  wire[63:0] T296;
  wire[63:0] scr_rdata_18;
  wire[63:0] scr_rdata_19;
  wire T297;
  wire T298;
  wire[63:0] T299;
  wire[63:0] T300;
  wire[63:0] scr_rdata_20;
  wire[63:0] scr_rdata_21;
  wire T301;
  wire[63:0] T302;
  wire[63:0] scr_rdata_22;
  wire[63:0] scr_rdata_23;
  wire T303;
  wire T304;
  wire T305;
  wire[63:0] T306;
  wire[63:0] T307;
  wire[63:0] T308;
  wire[63:0] scr_rdata_24;
  wire[63:0] scr_rdata_25;
  wire T309;
  wire[63:0] T310;
  wire[63:0] scr_rdata_26;
  wire[63:0] scr_rdata_27;
  wire T311;
  wire T312;
  wire[63:0] T313;
  wire[63:0] T314;
  wire[63:0] scr_rdata_28;
  wire[63:0] scr_rdata_29;
  wire T315;
  wire[63:0] T316;
  wire[63:0] scr_rdata_30;
  wire[63:0] scr_rdata_31;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire[63:0] T322;
  wire[63:0] T323;
  wire[63:0] T324;
  wire[63:0] T325;
  wire[63:0] T326;
  wire[63:0] scr_rdata_32;
  wire[63:0] scr_rdata_33;
  wire T327;
  wire[63:0] T328;
  wire[63:0] scr_rdata_34;
  wire[63:0] scr_rdata_35;
  wire T329;
  wire T330;
  wire[63:0] T331;
  wire[63:0] T332;
  wire[63:0] scr_rdata_36;
  wire[63:0] scr_rdata_37;
  wire T333;
  wire[63:0] T334;
  wire[63:0] scr_rdata_38;
  wire[63:0] scr_rdata_39;
  wire T335;
  wire T336;
  wire T337;
  wire[63:0] T338;
  wire[63:0] T339;
  wire[63:0] T340;
  wire[63:0] scr_rdata_40;
  wire[63:0] scr_rdata_41;
  wire T341;
  wire[63:0] T342;
  wire[63:0] scr_rdata_42;
  wire[63:0] scr_rdata_43;
  wire T343;
  wire T344;
  wire[63:0] T345;
  wire[63:0] T346;
  wire[63:0] scr_rdata_44;
  wire[63:0] scr_rdata_45;
  wire T347;
  wire[63:0] T348;
  wire[63:0] scr_rdata_46;
  wire[63:0] scr_rdata_47;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire[63:0] T353;
  wire[63:0] T354;
  wire[63:0] T355;
  wire[63:0] T356;
  wire[63:0] scr_rdata_48;
  wire[63:0] scr_rdata_49;
  wire T357;
  wire[63:0] T358;
  wire[63:0] scr_rdata_50;
  wire[63:0] scr_rdata_51;
  wire T359;
  wire T360;
  wire[63:0] T361;
  wire[63:0] T362;
  wire[63:0] scr_rdata_52;
  wire[63:0] scr_rdata_53;
  wire T363;
  wire[63:0] T364;
  wire[63:0] scr_rdata_54;
  wire[63:0] scr_rdata_55;
  wire T365;
  wire T366;
  wire T367;
  wire[63:0] T368;
  wire[63:0] T369;
  wire[63:0] T370;
  wire[63:0] scr_rdata_56;
  wire[63:0] scr_rdata_57;
  wire T371;
  wire[63:0] T372;
  wire[63:0] scr_rdata_58;
  wire[63:0] scr_rdata_59;
  wire T373;
  wire T374;
  wire[63:0] T375;
  wire[63:0] T376;
  wire[63:0] scr_rdata_60;
  wire[63:0] scr_rdata_61;
  wire T377;
  wire[63:0] T378;
  wire[63:0] scr_rdata_62;
  wire[63:0] scr_rdata_63;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[63:0] tx_header;
  wire[15:0] T388;
  wire[3:0] tx_cmd_ext;
  wire[2:0] tx_cmd;
  wire[47:0] T389;
  reg [7:0] seqno;
  wire[7:0] T390;
  wire[7:0] T391;
  wire T392;
  wire T393;
  wire T394;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    addr = {2{$random}};
    rx_shifter = {2{$random}};
    rx_count = {1{$random}};
    size = {1{$random}};
    cmd = {1{$random}};
    tx_count = {1{$random}};
    state = {1{$random}};
    mem_acked = {1{$random}};
    pos = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      packet_ram[initvar] = {2{$random}};
    mem_gxid = {1{$random}};
    mem_gsrc = {1{$random}};
    mem_needs_ack = {1{$random}};
    R231 = {1{$random}};
    R242 = {1{$random}};
    pcrReadData = {2{$random}};
    seqno = {1{$random}};
  end
`endif

  assign T0 = T1[2'h3:1'h0];
  assign T1 = T160 ? T146 : T2;
  assign T2 = {T10, T3};
  assign T3 = {T7, T4};
  assign T4 = {T6, T5};
  assign T5 = 4'h0;
  assign T6 = 3'h0;
  assign T7 = {T9, T8};
  assign T8 = 6'h0;
  assign T9 = 3'h2;
  assign T10 = {T14, T11};
  assign T11 = {T13, T12};
  assign T12 = 512'h0;
  assign T13 = 4'h0;
  assign T14 = T15;
  assign T15 = init_addr[5'h19:1'h0];
  assign init_addr = T16 >> 2'h3;
  assign T16 = addr;
  assign T17 = T127 ? T145 : T18;
  assign T18 = T23 ? T19 : addr;
  assign T19 = rx_shifter_in[6'h3f:5'h18];
  assign rx_shifter_in = {io_host_in_bits, T20};
  assign T20 = rx_shifter[6'h3f:5'h10];
  assign T21 = T22 ? rx_shifter_in : rx_shifter;
  assign T22 = io_host_in_valid & io_host_in_ready;
  assign T23 = T22 & T24;
  assign T24 = rx_count == 15'h3;
  assign T25 = reset ? 15'h0 : T26;
  assign T26 = T29 ? 15'h0 : T27;
  assign T27 = T22 ? T28 : rx_count;
  assign T28 = rx_count + 15'h1;
  assign T29 = T61 & T30;
  assign T30 = T55 == T31;
  assign T31 = {1'h0, tx_size};
  assign tx_size = T34 ? size : 12'h0;
  assign T32 = T23 ? T33 : size;
  assign T33 = rx_shifter_in[4'hf:3'h4];
  assign T34 = T42 & T35;
  assign T35 = T39 | T36;
  assign T36 = cmd == 4'h3;
  assign T37 = T23 ? T38 : cmd;
  assign T38 = rx_shifter_in[2'h3:1'h0];
  assign T39 = T41 | T40;
  assign T40 = cmd == 4'h2;
  assign T41 = cmd == 4'h0;
  assign T42 = nack ^ 1'h1;
  assign nack = T52 ? bad_mem_packet : T43;
  assign T43 = T45 ? T44 : 1'h1;
  assign T44 = size != 12'h1;
  assign T45 = T47 | T46;
  assign T46 = cmd == 4'h3;
  assign T47 = cmd == 4'h2;
  assign bad_mem_packet = T50 | T48;
  assign T48 = T49 != 3'h0;
  assign T49 = addr[2'h2:1'h0];
  assign T50 = T51 != 3'h0;
  assign T51 = size[2'h2:1'h0];
  assign T52 = T54 | T53;
  assign T53 = cmd == 4'h1;
  assign T54 = cmd == 4'h0;
  assign T55 = tx_count[4'he:2'h2];
  assign T56 = reset ? 15'h0 : T57;
  assign T57 = T29 ? 15'h0 : T58;
  assign T58 = T60 ? T59 : tx_count;
  assign T59 = tx_count + 15'h1;
  assign T60 = io_host_out_valid & io_host_out_ready;
  assign T61 = T72 & tx_done;
  assign tx_done = T69 & T62;
  assign T62 = T67 | T63;
  assign T63 = T66 & T64;
  assign T64 = packet_ram_raddr == 3'h7;
  assign packet_ram_raddr = T65 - 3'h1;
  assign T65 = T55[2'h2:1'h0];
  assign T66 = 13'h0 < T55;
  assign T67 = T55 == T68;
  assign T68 = {1'h0, tx_size};
  assign T69 = io_host_out_ready & T70;
  assign T70 = T71 == 2'h3;
  assign T71 = tx_count[1'h1:1'h0];
  assign T72 = state == 4'h8;
  assign T73 = reset ? 4'h0 : T74;
  assign T74 = T142 ? 4'h8 : T75;
  assign T75 = io_cpu_0_pcr_rep_valid ? 4'h8 : T76;
  assign T76 = T135 ? 4'h8 : T77;
  assign T77 = T134 ? 4'h2 : T78;
  assign T78 = T61 ? T130 : T79;
  assign T79 = T127 ? T120 : T80;
  assign T80 = T119 ? 4'h7 : T81;
  assign T81 = T112 ? 4'h7 : T82;
  assign T82 = T110 ? 4'h5 : T83;
  assign T83 = T108 ? 4'h6 : T84;
  assign T84 = T94 ? T85 : state;
  assign T85 = T93 ? 4'h3 : T86;
  assign T86 = T92 ? 4'h4 : T87;
  assign T87 = T88 ? 4'h1 : 4'h8;
  assign T88 = T91 | T89;
  assign T89 = rx_cmd == 4'h3;
  assign rx_cmd = T90 ? T38 : cmd;
  assign T90 = rx_word_count == 13'h0;
  assign rx_word_count = rx_count >> 2'h2;
  assign T91 = rx_cmd == 4'h2;
  assign T92 = rx_cmd == 4'h1;
  assign T93 = rx_cmd == 4'h0;
  assign T94 = T107 & rx_done;
  assign rx_done = rx_word_done & T95;
  assign T95 = T104 ? T101 : T96;
  assign T96 = T99 | T97;
  assign T97 = T98 == 3'h0;
  assign T98 = rx_word_count[2'h2:1'h0];
  assign T99 = rx_word_count == T100;
  assign T100 = {1'h0, size};
  assign T101 = T103 & T102;
  assign T102 = T38 != 4'h3;
  assign T103 = T38 != 4'h1;
  assign T104 = rx_word_count == 13'h0;
  assign rx_word_done = io_host_in_valid & T105;
  assign T105 = T106 == 2'h3;
  assign T106 = rx_count[1'h1:1'h0];
  assign T107 = state == 4'h0;
  assign T108 = T109 & acq_q_io_enq_ready;
  assign T109 = state == 4'h4;
  assign T110 = T111 & acq_q_io_enq_ready;
  assign T111 = state == 4'h3;
  assign T112 = T118 & mem_acked;
  assign T113 = reset ? 1'h0 : T114;
  assign T114 = T117 ? 1'h0 : T115;
  assign T115 = T112 ? 1'h0 : T116;
  assign T116 = io_mem_grant_valid ? 1'h1 : mem_acked;
  assign T117 = state == 4'h5;
  assign T118 = state == 4'h6;
  assign T119 = T117 & io_mem_grant_valid;
  assign T120 = T121 ? 4'h8 : 4'h0;
  assign T121 = T129 | T122;
  assign T122 = pos == 9'h1;
  assign T123 = T127 ? T126 : T124;
  assign T124 = T23 ? T125 : pos;
  assign T125 = rx_shifter_in[4'hf:3'h7];
  assign T126 = pos - 9'h1;
  assign T127 = T128 & io_mem_finish_ready;
  assign T128 = state == 4'h7;
  assign T129 = cmd == 4'h0;
  assign T130 = T131 ? 4'h3 : 4'h0;
  assign T131 = T133 & T132;
  assign T132 = pos != 9'h0;
  assign T133 = cmd == 4'h0;
  assign T134 = io_cpu_0_pcr_req_valid & io_cpu_0_pcr_req_ready;
  assign T135 = T138 & T136;
  assign T136 = T137 == 5'h1d;
  assign T137 = addr[3'h4:1'h0];
  assign T138 = T141 & T139;
  assign T139 = T140 == 2'h0;
  assign T140 = addr[5'h15:5'h14];
  assign T141 = state == 4'h1;
  assign T142 = T144 & T143;
  assign T143 = T140 == 2'h3;
  assign T144 = state == 4'h1;
  assign T145 = addr + 40'h8;
  assign T146 = {T154, T147};
  assign T147 = {T151, T148};
  assign T148 = {T150, T149};
  assign T149 = 4'h0;
  assign T150 = 3'h0;
  assign T151 = {T153, T152};
  assign T152 = 6'h0;
  assign T153 = 3'h3;
  assign T154 = {T158, T155};
  assign T155 = {T157, T156};
  assign T156 = 512'h0;
  assign T157 = 4'h0;
  assign T158 = T159;
  assign T159 = init_addr[5'h19:1'h0];
  assign T160 = cmd == 4'h1;
  assign T161 = T1[3'h6:3'h4];
  assign T162 = T1[4'hc:3'h7];
  assign T163 = T1[4'hf:4'hd];
  assign T164 = T1[10'h20f:5'h10];
  assign T165 = T1[10'h213:10'h210];
  assign T166 = T1[10'h22d:10'h214];
  assign T167 = T169 | T168;
  assign T168 = state == 4'h4;
  assign T169 = state == 4'h3;
  assign io_scr_wdata = T170;
  assign T170 = packet_ram_0[3'h0] ^ packet_ram_1[3'h0] ^ packet_ram_2[3'h0] ^ packet_ram_3[3'h0] ^ packet_ram_4[3'h0] ^ packet_ram_5[3'h0] ^ packet_ram_6[3'h0] ^ packet_ram_7[3'h0] ^ packet_ram_8[3'h0];
  wire [63:0] packet_ram_w8 = packet_ram_0[3'h7] ^ packet_ram_1[3'h7] ^ packet_ram_2[3'h7] ^ packet_ram_3[3'h7] ^ packet_ram_4[3'h7] ^ packet_ram_5[3'h7] ^ packet_ram_6[3'h7] ^ packet_ram_7[3'h7];
  always @(posedge clk)
    if (T173)
      packet_ram_8[3'h7] <= T172 ^ packet_ram_w8;
  assign T172 = io_mem_grant_bits_payload_data[9'h1ff:9'h1c0];
  assign T173 = T174 & io_mem_grant_valid;
  assign T174 = state == 4'h5;
  wire [63:0] packet_ram_w7 = packet_ram_0[3'h6] ^ packet_ram_1[3'h6] ^ packet_ram_2[3'h6] ^ packet_ram_3[3'h6] ^ packet_ram_4[3'h6] ^ packet_ram_5[3'h6] ^ packet_ram_6[3'h6] ^ packet_ram_8[3'h6];
  always @(posedge clk)
    if (T177)
      packet_ram_7[3'h6] <= T176 ^ packet_ram_w7;
  assign T176 = io_mem_grant_bits_payload_data[9'h1bf:9'h180];
  assign T177 = T178 & io_mem_grant_valid;
  assign T178 = state == 4'h5;
  wire [63:0] packet_ram_w6 = packet_ram_0[3'h5] ^ packet_ram_1[3'h5] ^ packet_ram_2[3'h5] ^ packet_ram_3[3'h5] ^ packet_ram_4[3'h5] ^ packet_ram_5[3'h5] ^ packet_ram_7[3'h5] ^ packet_ram_8[3'h5];
  always @(posedge clk)
    if (T181)
      packet_ram_6[3'h5] <= T180 ^ packet_ram_w6;
  assign T180 = io_mem_grant_bits_payload_data[9'h17f:9'h140];
  assign T181 = T182 & io_mem_grant_valid;
  assign T182 = state == 4'h5;
  wire [63:0] packet_ram_w5 = packet_ram_0[3'h4] ^ packet_ram_1[3'h4] ^ packet_ram_2[3'h4] ^ packet_ram_3[3'h4] ^ packet_ram_4[3'h4] ^ packet_ram_6[3'h4] ^ packet_ram_7[3'h4] ^ packet_ram_8[3'h4];
  always @(posedge clk)
    if (T185)
      packet_ram_5[3'h4] <= T184 ^ packet_ram_w5;
  assign T184 = io_mem_grant_bits_payload_data[9'h13f:9'h100];
  assign T185 = T186 & io_mem_grant_valid;
  assign T186 = state == 4'h5;
  wire [63:0] packet_ram_w4 = packet_ram_0[3'h3] ^ packet_ram_1[3'h3] ^ packet_ram_2[3'h3] ^ packet_ram_3[3'h3] ^ packet_ram_5[3'h3] ^ packet_ram_6[3'h3] ^ packet_ram_7[3'h3] ^ packet_ram_8[3'h3];
  always @(posedge clk)
    if (T189)
      packet_ram_4[3'h3] <= T188 ^ packet_ram_w4;
  assign T188 = io_mem_grant_bits_payload_data[8'hff:8'hc0];
  assign T189 = T190 & io_mem_grant_valid;
  assign T190 = state == 4'h5;
  wire [63:0] packet_ram_w3 = packet_ram_0[3'h2] ^ packet_ram_1[3'h2] ^ packet_ram_2[3'h2] ^ packet_ram_4[3'h2] ^ packet_ram_5[3'h2] ^ packet_ram_6[3'h2] ^ packet_ram_7[3'h2] ^ packet_ram_8[3'h2];
  always @(posedge clk)
    if (T193)
      packet_ram_3[3'h2] <= T192 ^ packet_ram_w3;
  assign T192 = io_mem_grant_bits_payload_data[8'hbf:8'h80];
  assign T193 = T194 & io_mem_grant_valid;
  assign T194 = state == 4'h5;
  wire [63:0] packet_ram_w2 = packet_ram_0[3'h1] ^ packet_ram_1[3'h1] ^ packet_ram_3[3'h1] ^ packet_ram_4[3'h1] ^ packet_ram_5[3'h1] ^ packet_ram_6[3'h1] ^ packet_ram_7[3'h1] ^ packet_ram_8[3'h1];
  always @(posedge clk)
    if (T197)
      packet_ram_2[3'h1] <= T196 ^ packet_ram_w2;
  assign T196 = io_mem_grant_bits_payload_data[7'h7f:7'h40];
  assign T197 = T198 & io_mem_grant_valid;
  assign T198 = state == 4'h5;
  wire [63:0] packet_ram_w1 = packet_ram_0[3'h0] ^ packet_ram_2[3'h0] ^ packet_ram_3[3'h0] ^ packet_ram_4[3'h0] ^ packet_ram_5[3'h0] ^ packet_ram_6[3'h0] ^ packet_ram_7[3'h0] ^ packet_ram_8[3'h0];
  always @(posedge clk)
    if (T201)
      packet_ram_1[3'h0] <= T200 ^ packet_ram_w1;
  assign T200 = io_mem_grant_bits_payload_data[6'h3f:1'h0];
  assign T201 = T202 & io_mem_grant_valid;
  assign T202 = state == 4'h5;
  wire [63:0] packet_ram_w0 = packet_ram_1[T205] ^ packet_ram_2[T205] ^ packet_ram_3[T205] ^ packet_ram_4[T205] ^ packet_ram_5[T205] ^ packet_ram_6[T205] ^ packet_ram_7[T205] ^ packet_ram_8[T205];
  always @(posedge clk)
    if (T204)
      packet_ram_0[T205] <= rx_shifter_in ^ packet_ram_w0;
  assign T204 = rx_word_done & io_host_in_ready;
  assign T205 = T206 - 3'h1;
  assign T206 = rx_word_count[2'h2:1'h0];
  assign io_scr_waddr = T207;
  assign T207 = T208;
  assign T208 = addr[3'h5:1'h0];
  assign io_scr_wen = T209;
  assign T209 = T142 ? T210 : 1'h0;
  assign T210 = cmd == 4'h3;
  assign io_mem_release_valid = 1'h0;
  assign io_mem_probe_ready = 1'h0;
  assign io_mem_finish_bits_payload_master_xact_id = mem_gxid;
  assign T211 = io_mem_grant_valid ? io_mem_grant_bits_payload_master_xact_id : mem_gxid;
  assign io_mem_finish_bits_header_dst = mem_gsrc;
  assign T212 = io_mem_grant_valid ? io_mem_grant_bits_header_src : mem_gsrc;
  assign io_mem_finish_valid = T213;
  assign T213 = T216 & mem_needs_ack;
  assign T214 = io_mem_grant_valid ? T215 : mem_needs_ack;
  assign T215 = io_mem_grant_bits_payload_g_type != 4'h0;
  assign T216 = state == 4'h7;
  assign io_mem_grant_ready = 1'h1;
  assign io_mem_acquire_bits_payload_atomic_opcode = acq_q_io_deq_bits_atomic_opcode;
  assign io_mem_acquire_bits_payload_subword_addr = acq_q_io_deq_bits_subword_addr;
  assign io_mem_acquire_bits_payload_write_mask = acq_q_io_deq_bits_write_mask;
  assign io_mem_acquire_bits_payload_a_type = acq_q_io_deq_bits_a_type;
  assign io_mem_acquire_bits_payload_data = mem_req_data;
  assign mem_req_data = {T230, T217};
  assign T217 = {T229, T218};
  assign T218 = {T228, T219};
  assign T219 = {T227, T220};
  assign T220 = {T226, T221};
  assign T221 = {T225, T222};
  assign T222 = {T224, T223};
  assign T223 = packet_ram_0[3'h0] ^ packet_ram_1[3'h0] ^ packet_ram_2[3'h0] ^ packet_ram_3[3'h0] ^ packet_ram_4[3'h0] ^ packet_ram_5[3'h0] ^ packet_ram_6[3'h0] ^ packet_ram_7[3'h0] ^ packet_ram_8[3'h0];
  assign T224 = packet_ram_0[3'h1] ^ packet_ram_1[3'h1] ^ packet_ram_2[3'h1] ^ packet_ram_3[3'h1] ^ packet_ram_4[3'h1] ^ packet_ram_5[3'h1] ^ packet_ram_6[3'h1] ^ packet_ram_7[3'h1] ^ packet_ram_8[3'h1];
  assign T225 = packet_ram_0[3'h2] ^ packet_ram_1[3'h2] ^ packet_ram_2[3'h2] ^ packet_ram_3[3'h2] ^ packet_ram_4[3'h2] ^ packet_ram_5[3'h2] ^ packet_ram_6[3'h2] ^ packet_ram_7[3'h2] ^ packet_ram_8[3'h2];
  assign T226 = packet_ram_0[3'h3] ^ packet_ram_1[3'h3] ^ packet_ram_2[3'h3] ^ packet_ram_3[3'h3] ^ packet_ram_4[3'h3] ^ packet_ram_5[3'h3] ^ packet_ram_6[3'h3] ^ packet_ram_7[3'h3] ^ packet_ram_8[3'h3];
  assign T227 = packet_ram_0[3'h4] ^ packet_ram_1[3'h4] ^ packet_ram_2[3'h4] ^ packet_ram_3[3'h4] ^ packet_ram_4[3'h4] ^ packet_ram_5[3'h4] ^ packet_ram_6[3'h4] ^ packet_ram_7[3'h4] ^ packet_ram_8[3'h4];
  assign T228 = packet_ram_0[3'h5] ^ packet_ram_1[3'h5] ^ packet_ram_2[3'h5] ^ packet_ram_3[3'h5] ^ packet_ram_4[3'h5] ^ packet_ram_5[3'h5] ^ packet_ram_6[3'h5] ^ packet_ram_7[3'h5] ^ packet_ram_8[3'h5];
  assign T229 = packet_ram_0[3'h6] ^ packet_ram_1[3'h6] ^ packet_ram_2[3'h6] ^ packet_ram_3[3'h6] ^ packet_ram_4[3'h6] ^ packet_ram_5[3'h6] ^ packet_ram_6[3'h6] ^ packet_ram_7[3'h6] ^ packet_ram_8[3'h6];
  assign T230 = packet_ram_0[3'h7] ^ packet_ram_1[3'h7] ^ packet_ram_2[3'h7] ^ packet_ram_3[3'h7] ^ packet_ram_4[3'h7] ^ packet_ram_5[3'h7] ^ packet_ram_6[3'h7] ^ packet_ram_7[3'h7] ^ packet_ram_8[3'h7];
  assign io_mem_acquire_bits_payload_client_xact_id = acq_q_io_deq_bits_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = acq_q_io_deq_bits_addr;
  assign io_mem_acquire_bits_header_dst = 2'h0;
  assign io_mem_acquire_bits_header_src = 2'h2;
  assign io_mem_acquire_valid = acq_q_io_deq_valid;
  assign io_cpu_0_ipi_rep_valid = R231;
  assign T232 = reset ? 1'h0 : T233;
  assign T233 = T235 ? 1'h1 : T234;
  assign T234 = io_cpu_0_ipi_rep_ready ? 1'h0 : R231;
  assign T235 = io_cpu_0_ipi_req_valid & T236;
  assign T236 = io_cpu_0_ipi_req_bits == 1'h0;
  assign io_cpu_0_ipi_req_ready = 1'h1;
  assign io_cpu_0_pcr_rep_ready = 1'h1;
  assign io_cpu_0_pcr_req_bits_data = T170;
  assign io_cpu_0_pcr_req_bits_addr = T137;
  assign io_cpu_0_pcr_req_bits_rw = T237;
  assign T237 = cmd == 4'h3;
  assign io_cpu_0_pcr_req_valid = T238;
  assign T238 = T240 & T239;
  assign T239 = T137 != 5'h1d;
  assign T240 = T241 & T139;
  assign T241 = state == 4'h1;
  assign io_cpu_0_reset = R242;
  assign T243 = reset ? 1'h1 : T244;
  assign T244 = T246 ? T245 : R242;
  assign T245 = T170[1'h0:1'h0];
  assign T246 = T135 & T247;
  assign T247 = cmd == 4'h3;
  assign io_host_debug_stats_pcr = io_cpu_0_debug_stats_pcr;
  assign io_host_out_bits = T248;
  assign T248 = T249[4'hf:1'h0];
  assign T249 = tx_data >> T250;
  assign T250 = {T251, 4'h0};
  assign T251 = tx_count[1'h1:1'h0];
  assign tx_data = T392 ? tx_header : T252;
  assign T252 = T385 ? pcrReadData : T253;
  assign T253 = packet_ram_0[packet_ram_raddr] ^ packet_ram_1[packet_ram_raddr] ^ packet_ram_2[packet_ram_raddr] ^ packet_ram_3[packet_ram_raddr] ^ packet_ram_4[packet_ram_raddr] ^ packet_ram_5[packet_ram_raddr] ^ packet_ram_6[packet_ram_raddr] ^ packet_ram_7[packet_ram_raddr] ^ packet_ram_8[packet_ram_raddr];
  assign T254 = T142 ? T258 : T255;
  assign T255 = io_cpu_0_pcr_rep_valid ? io_cpu_0_pcr_rep_bits : T256;
  assign T256 = T135 ? T257 : pcrReadData;
  assign T257 = {63'h0, R242};
  assign T258 = T384 ? T322 : T259;
  assign T259 = T321 ? T291 : T260;
  assign T260 = T290 ? T276 : T261;
  assign T261 = T275 ? T269 : T262;
  assign T262 = T268 ? T266 : T263;
  assign T263 = T264 ? scr_rdata_1 : scr_rdata_0;
  assign scr_rdata_0 = 64'h1;
  assign scr_rdata_1 = 64'h1000;
  assign T264 = T265[1'h0:1'h0];
  assign T265 = T208;
  assign T266 = T267 ? scr_rdata_3 : scr_rdata_2;
  assign scr_rdata_2 = io_scr_rdata_2;
  assign scr_rdata_3 = io_scr_rdata_3;
  assign T267 = T265[1'h0:1'h0];
  assign T268 = T265[1'h1:1'h1];
  assign T269 = T274 ? T272 : T270;
  assign T270 = T271 ? scr_rdata_5 : scr_rdata_4;
  assign scr_rdata_4 = io_scr_rdata_4;
  assign scr_rdata_5 = io_scr_rdata_5;
  assign T271 = T265[1'h0:1'h0];
  assign T272 = T273 ? scr_rdata_7 : scr_rdata_6;
  assign scr_rdata_6 = io_scr_rdata_6;
  assign scr_rdata_7 = io_scr_rdata_7;
  assign T273 = T265[1'h0:1'h0];
  assign T274 = T265[1'h1:1'h1];
  assign T275 = T265[2'h2:2'h2];
  assign T276 = T289 ? T283 : T277;
  assign T277 = T282 ? T280 : T278;
  assign T278 = T279 ? scr_rdata_9 : scr_rdata_8;
  assign scr_rdata_8 = io_scr_rdata_8;
  assign scr_rdata_9 = io_scr_rdata_9;
  assign T279 = T265[1'h0:1'h0];
  assign T280 = T281 ? scr_rdata_11 : scr_rdata_10;
  assign scr_rdata_10 = io_scr_rdata_10;
  assign scr_rdata_11 = io_scr_rdata_11;
  assign T281 = T265[1'h0:1'h0];
  assign T282 = T265[1'h1:1'h1];
  assign T283 = T288 ? T286 : T284;
  assign T284 = T285 ? scr_rdata_13 : scr_rdata_12;
  assign scr_rdata_12 = io_scr_rdata_12;
  assign scr_rdata_13 = io_scr_rdata_13;
  assign T285 = T265[1'h0:1'h0];
  assign T286 = T287 ? scr_rdata_15 : scr_rdata_14;
  assign scr_rdata_14 = io_scr_rdata_14;
  assign scr_rdata_15 = io_scr_rdata_15;
  assign T287 = T265[1'h0:1'h0];
  assign T288 = T265[1'h1:1'h1];
  assign T289 = T265[2'h2:2'h2];
  assign T290 = T265[2'h3:2'h3];
  assign T291 = T320 ? T306 : T292;
  assign T292 = T305 ? T299 : T293;
  assign T293 = T298 ? T296 : T294;
  assign T294 = T295 ? scr_rdata_17 : scr_rdata_16;
  assign scr_rdata_16 = io_scr_rdata_16;
  assign scr_rdata_17 = io_scr_rdata_17;
  assign T295 = T265[1'h0:1'h0];
  assign T296 = T297 ? scr_rdata_19 : scr_rdata_18;
  assign scr_rdata_18 = io_scr_rdata_18;
  assign scr_rdata_19 = io_scr_rdata_19;
  assign T297 = T265[1'h0:1'h0];
  assign T298 = T265[1'h1:1'h1];
  assign T299 = T304 ? T302 : T300;
  assign T300 = T301 ? scr_rdata_21 : scr_rdata_20;
  assign scr_rdata_20 = io_scr_rdata_20;
  assign scr_rdata_21 = io_scr_rdata_21;
  assign T301 = T265[1'h0:1'h0];
  assign T302 = T303 ? scr_rdata_23 : scr_rdata_22;
  assign scr_rdata_22 = io_scr_rdata_22;
  assign scr_rdata_23 = io_scr_rdata_23;
  assign T303 = T265[1'h0:1'h0];
  assign T304 = T265[1'h1:1'h1];
  assign T305 = T265[2'h2:2'h2];
  assign T306 = T319 ? T313 : T307;
  assign T307 = T312 ? T310 : T308;
  assign T308 = T309 ? scr_rdata_25 : scr_rdata_24;
  assign scr_rdata_24 = io_scr_rdata_24;
  assign scr_rdata_25 = io_scr_rdata_25;
  assign T309 = T265[1'h0:1'h0];
  assign T310 = T311 ? scr_rdata_27 : scr_rdata_26;
  assign scr_rdata_26 = io_scr_rdata_26;
  assign scr_rdata_27 = io_scr_rdata_27;
  assign T311 = T265[1'h0:1'h0];
  assign T312 = T265[1'h1:1'h1];
  assign T313 = T318 ? T316 : T314;
  assign T314 = T315 ? scr_rdata_29 : scr_rdata_28;
  assign scr_rdata_28 = io_scr_rdata_28;
  assign scr_rdata_29 = io_scr_rdata_29;
  assign T315 = T265[1'h0:1'h0];
  assign T316 = T317 ? scr_rdata_31 : scr_rdata_30;
  assign scr_rdata_30 = io_scr_rdata_30;
  assign scr_rdata_31 = io_scr_rdata_31;
  assign T317 = T265[1'h0:1'h0];
  assign T318 = T265[1'h1:1'h1];
  assign T319 = T265[2'h2:2'h2];
  assign T320 = T265[2'h3:2'h3];
  assign T321 = T265[3'h4:3'h4];
  assign T322 = T383 ? T353 : T323;
  assign T323 = T352 ? T338 : T324;
  assign T324 = T337 ? T331 : T325;
  assign T325 = T330 ? T328 : T326;
  assign T326 = T327 ? scr_rdata_33 : scr_rdata_32;
  assign scr_rdata_32 = io_scr_rdata_32;
  assign scr_rdata_33 = io_scr_rdata_33;
  assign T327 = T265[1'h0:1'h0];
  assign T328 = T329 ? scr_rdata_35 : scr_rdata_34;
  assign scr_rdata_34 = io_scr_rdata_34;
  assign scr_rdata_35 = io_scr_rdata_35;
  assign T329 = T265[1'h0:1'h0];
  assign T330 = T265[1'h1:1'h1];
  assign T331 = T336 ? T334 : T332;
  assign T332 = T333 ? scr_rdata_37 : scr_rdata_36;
  assign scr_rdata_36 = io_scr_rdata_36;
  assign scr_rdata_37 = io_scr_rdata_37;
  assign T333 = T265[1'h0:1'h0];
  assign T334 = T335 ? scr_rdata_39 : scr_rdata_38;
  assign scr_rdata_38 = io_scr_rdata_38;
  assign scr_rdata_39 = io_scr_rdata_39;
  assign T335 = T265[1'h0:1'h0];
  assign T336 = T265[1'h1:1'h1];
  assign T337 = T265[2'h2:2'h2];
  assign T338 = T351 ? T345 : T339;
  assign T339 = T344 ? T342 : T340;
  assign T340 = T341 ? scr_rdata_41 : scr_rdata_40;
  assign scr_rdata_40 = io_scr_rdata_40;
  assign scr_rdata_41 = io_scr_rdata_41;
  assign T341 = T265[1'h0:1'h0];
  assign T342 = T343 ? scr_rdata_43 : scr_rdata_42;
  assign scr_rdata_42 = io_scr_rdata_42;
  assign scr_rdata_43 = io_scr_rdata_43;
  assign T343 = T265[1'h0:1'h0];
  assign T344 = T265[1'h1:1'h1];
  assign T345 = T350 ? T348 : T346;
  assign T346 = T347 ? scr_rdata_45 : scr_rdata_44;
  assign scr_rdata_44 = io_scr_rdata_44;
  assign scr_rdata_45 = io_scr_rdata_45;
  assign T347 = T265[1'h0:1'h0];
  assign T348 = T349 ? scr_rdata_47 : scr_rdata_46;
  assign scr_rdata_46 = io_scr_rdata_46;
  assign scr_rdata_47 = io_scr_rdata_47;
  assign T349 = T265[1'h0:1'h0];
  assign T350 = T265[1'h1:1'h1];
  assign T351 = T265[2'h2:2'h2];
  assign T352 = T265[2'h3:2'h3];
  assign T353 = T382 ? T368 : T354;
  assign T354 = T367 ? T361 : T355;
  assign T355 = T360 ? T358 : T356;
  assign T356 = T357 ? scr_rdata_49 : scr_rdata_48;
  assign scr_rdata_48 = io_scr_rdata_48;
  assign scr_rdata_49 = io_scr_rdata_49;
  assign T357 = T265[1'h0:1'h0];
  assign T358 = T359 ? scr_rdata_51 : scr_rdata_50;
  assign scr_rdata_50 = io_scr_rdata_50;
  assign scr_rdata_51 = io_scr_rdata_51;
  assign T359 = T265[1'h0:1'h0];
  assign T360 = T265[1'h1:1'h1];
  assign T361 = T366 ? T364 : T362;
  assign T362 = T363 ? scr_rdata_53 : scr_rdata_52;
  assign scr_rdata_52 = io_scr_rdata_52;
  assign scr_rdata_53 = io_scr_rdata_53;
  assign T363 = T265[1'h0:1'h0];
  assign T364 = T365 ? scr_rdata_55 : scr_rdata_54;
  assign scr_rdata_54 = io_scr_rdata_54;
  assign scr_rdata_55 = io_scr_rdata_55;
  assign T365 = T265[1'h0:1'h0];
  assign T366 = T265[1'h1:1'h1];
  assign T367 = T265[2'h2:2'h2];
  assign T368 = T381 ? T375 : T369;
  assign T369 = T374 ? T372 : T370;
  assign T370 = T371 ? scr_rdata_57 : scr_rdata_56;
  assign scr_rdata_56 = io_scr_rdata_56;
  assign scr_rdata_57 = io_scr_rdata_57;
  assign T371 = T265[1'h0:1'h0];
  assign T372 = T373 ? scr_rdata_59 : scr_rdata_58;
  assign scr_rdata_58 = io_scr_rdata_58;
  assign scr_rdata_59 = io_scr_rdata_59;
  assign T373 = T265[1'h0:1'h0];
  assign T374 = T265[1'h1:1'h1];
  assign T375 = T380 ? T378 : T376;
  assign T376 = T377 ? scr_rdata_61 : scr_rdata_60;
  assign scr_rdata_60 = io_scr_rdata_60;
  assign scr_rdata_61 = io_scr_rdata_61;
  assign T377 = T265[1'h0:1'h0];
  assign T378 = T379 ? scr_rdata_63 : scr_rdata_62;
  assign scr_rdata_62 = io_scr_rdata_62;
  assign scr_rdata_63 = io_scr_rdata_63;
  assign T379 = T265[1'h0:1'h0];
  assign T380 = T265[1'h1:1'h1];
  assign T381 = T265[2'h2:2'h2];
  assign T382 = T265[2'h3:2'h3];
  assign T383 = T265[3'h4:3'h4];
  assign T384 = T265[3'h5:3'h5];
  assign T385 = T387 | T386;
  assign T386 = cmd == 4'h3;
  assign T387 = cmd == 4'h2;
  assign tx_header = {T389, T388};
  assign T388 = {tx_size, tx_cmd_ext};
  assign tx_cmd_ext = {1'h0, tx_cmd};
  assign tx_cmd = nack ? 3'h5 : 3'h4;
  assign T389 = {addr, seqno};
  assign T390 = T23 ? T391 : seqno;
  assign T391 = rx_shifter_in[5'h17:5'h10];
  assign T392 = T55 == 13'h0;
  assign io_host_out_valid = T393;
  assign T393 = state == 4'h8;
  assign io_host_in_ready = T394;
  assign T394 = state == 4'h0;
  Queue_2 acq_q(.clk(clk), .reset(reset),
       .io_enq_ready( acq_q_io_enq_ready ),
       .io_enq_valid( T167 ),
       .io_enq_bits_addr( T166 ),
       .io_enq_bits_client_xact_id( T165 ),
       .io_enq_bits_data( T164 ),
       .io_enq_bits_a_type( T163 ),
       .io_enq_bits_write_mask( T162 ),
       .io_enq_bits_subword_addr( T161 ),
       .io_enq_bits_atomic_opcode( T0 ),
       .io_deq_ready( io_mem_acquire_ready ),
       .io_deq_valid( acq_q_io_deq_valid ),
       .io_deq_bits_addr( acq_q_io_deq_bits_addr ),
       .io_deq_bits_client_xact_id( acq_q_io_deq_bits_client_xact_id ),
       //.io_deq_bits_data(  )
       .io_deq_bits_a_type( acq_q_io_deq_bits_a_type ),
       .io_deq_bits_write_mask( acq_q_io_deq_bits_write_mask ),
       .io_deq_bits_subword_addr( acq_q_io_deq_bits_subword_addr ),
       .io_deq_bits_atomic_opcode( acq_q_io_deq_bits_atomic_opcode )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(T127) begin
      addr <= T145;
    end else if(T23) begin
      addr <= T19;
    end
    if(T22) begin
      rx_shifter <= rx_shifter_in;
    end
    if(reset) begin
      rx_count <= 15'h0;
    end else if(T29) begin
      rx_count <= 15'h0;
    end else if(T22) begin
      rx_count <= T28;
    end
    if(T23) begin
      size <= T33;
    end
    if(T23) begin
      cmd <= T38;
    end
    if(reset) begin
      tx_count <= 15'h0;
    end else if(T29) begin
      tx_count <= 15'h0;
    end else if(T60) begin
      tx_count <= T59;
    end
    if(reset) begin
      state <= 4'h0;
    end else if(T142) begin
      state <= 4'h8;
    end else if(io_cpu_0_pcr_rep_valid) begin
      state <= 4'h8;
    end else if(T135) begin
      state <= 4'h8;
    end else if(T134) begin
      state <= 4'h2;
    end else if(T61) begin
      state <= T130;
    end else if(T127) begin
      state <= T120;
    end else if(T119) begin
      state <= 4'h7;
    end else if(T112) begin
      state <= 4'h7;
    end else if(T110) begin
      state <= 4'h5;
    end else if(T108) begin
      state <= 4'h6;
    end else if(T94) begin
      state <= T85;
    end
    if(reset) begin
      mem_acked <= 1'h0;
    end else if(T117) begin
      mem_acked <= 1'h0;
    end else if(T112) begin
      mem_acked <= 1'h0;
    end else if(io_mem_grant_valid) begin
      mem_acked <= 1'h1;
    end
    if(T127) begin
      pos <= T126;
    end else if(T23) begin
      pos <= T125;
    end
    if(io_mem_grant_valid) begin
      mem_gxid <= io_mem_grant_bits_payload_master_xact_id;
    end
    if(io_mem_grant_valid) begin
      mem_gsrc <= io_mem_grant_bits_header_src;
    end
    if(io_mem_grant_valid) begin
      mem_needs_ack <= T215;
    end
    if(reset) begin
      R231 <= 1'h0;
    end else if(T235) begin
      R231 <= 1'h1;
    end else if(io_cpu_0_ipi_rep_ready) begin
      R231 <= 1'h0;
    end
    if(reset) begin
      R242 <= 1'h1;
    end else if(T246) begin
      R242 <= T245;
    end
    if(T142) begin
      pcrReadData <= T258;
    end else if(io_cpu_0_pcr_rep_valid) begin
      pcrReadData <= io_cpu_0_pcr_rep_bits;
    end else if(T135) begin
      pcrReadData <= T257;
    end
    if(T23) begin
      seqno <= T391;
    end
  end
endmodule

module VoluntaryReleaseTracker(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [3:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[3:0] io_inner_grant_bits_payload_client_xact_id,
    output[3:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [3:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    //output[1:0] io_inner_probe_bits_header_src
    //output[1:0] io_inner_probe_bits_header_dst
    //output[25:0] io_inner_probe_bits_payload_addr
    //output[3:0] io_inner_probe_bits_payload_master_xact_id
    //output[1:0] io_inner_probe_bits_payload_p_type
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [3:0] io_inner_release_bits_payload_client_xact_id,
    input [3:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[3:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [3:0] io_outer_grant_bits_payload_client_xact_id,
    input [3:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[3:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [1:0] state;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  reg [25:0] xact_addr;
  wire[25:0] T21;
  wire[3:0] T22;
  wire[2:0] T23;
  wire[5:0] T24;
  wire[2:0] T25;
  wire[511:0] T26;
  reg [511:0] xact_data;
  wire[511:0] T27;
  wire[3:0] T28;
  wire[25:0] T29;
  wire[3:0] T30;
  wire[3:0] T31;
  wire T32;
  reg [2:0] xact_r_type;
  wire[2:0] T33;
  wire[3:0] T34;
  wire[3:0] T35;
  reg [3:0] xact_client_xact_id;
  wire[3:0] T36;
  wire[511:0] T37;
  wire[1:0] T38;
  reg  init_client_id;
  wire T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire[1:0] T42;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    xact_r_type = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T20 & T1;
  assign T1 = state != 2'h0;
  assign T2 = reset ? 2'h0 : T3;
  assign T3 = T18 ? 2'h0 : T4;
  assign T4 = T16 ? 2'h2 : T5;
  assign T5 = T14 ? T6 : state;
  assign T6 = T7 ? 2'h1 : 2'h2;
  assign T7 = T9 | T8;
  assign T8 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T9 = T11 | T10;
  assign T10 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T11 = T13 | T12;
  assign T12 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T13 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T14 = T15 & io_inner_release_valid;
  assign T15 = 2'h0 == state;
  assign T16 = T17 & io_outer_acquire_ready;
  assign T17 = 2'h1 == state;
  assign T18 = T19 & io_inner_grant_ready;
  assign T19 = 2'h2 == state;
  assign T20 = xact_addr == io_inner_release_bits_payload_addr;
  assign T21 = T14 ? io_inner_release_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = 1'h0;
  assign io_outer_grant_ready = 1'h0;
  assign io_outer_acquire_bits_payload_atomic_opcode = T22;
  assign T22 = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T23;
  assign T23 = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T24;
  assign T24 = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T25;
  assign T25 = 3'h3;
  assign io_outer_acquire_bits_payload_data = T26;
  assign T26 = xact_data;
  assign T27 = T14 ? io_inner_release_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T28;
  assign T28 = 4'h0;
  assign io_outer_acquire_bits_payload_addr = T29;
  assign T29 = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T17;
  assign io_inner_release_ready = T15;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_grant_bits_payload_g_type = T30;
  assign T30 = T31;
  assign T31 = T32 ? 4'h0 : 4'h3;
  assign T32 = xact_r_type == 3'h0;
  assign T33 = T14 ? io_inner_release_bits_payload_r_type : xact_r_type;
  assign io_inner_grant_bits_payload_master_xact_id = T34;
  assign T34 = 4'h0;
  assign io_inner_grant_bits_payload_client_xact_id = T35;
  assign T35 = xact_client_xact_id;
  assign T36 = T14 ? io_inner_release_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T37;
  assign T37 = 512'h0;
  assign io_inner_grant_bits_header_dst = T38;
  assign T38 = {1'h0, init_client_id};
  assign T39 = T40[1'h0:1'h0];
  assign T40 = reset ? 2'h0 : T41;
  assign T41 = T14 ? io_inner_release_bits_header_src : T42;
  assign T42 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T19;
  assign io_inner_acquire_ready = 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else if(T18) begin
      state <= 2'h0;
    end else if(T16) begin
      state <= 2'h2;
    end else if(T14) begin
      state <= T6;
    end
    if(T14) begin
      xact_addr <= io_inner_release_bits_payload_addr;
    end
    if(T14) begin
      xact_data <= io_inner_release_bits_payload_data;
    end
    if(T14) begin
      xact_r_type <= io_inner_release_bits_payload_r_type;
    end
    if(T14) begin
      xact_client_xact_id <= io_inner_release_bits_payload_client_xact_id;
    end
    init_client_id <= T39;
  end
endmodule

module AcquireTracker_0(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [3:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[3:0] io_inner_grant_bits_payload_client_xact_id,
    output[3:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [3:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[3:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [3:0] io_inner_release_bits_payload_client_xact_id,
    input [3:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[3:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [3:0] io_outer_grant_bits_payload_client_xact_id,
    input [3:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[3:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] probe_initial_flags;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  reg [2:0] xact_a_type;
  wire[2:0] T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  reg  release_count;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[2:0] T62;
  wire[2:0] T63;
  wire T64;
  wire T65;
  wire[2:0] T66;
  wire T67;
  wire[3:0] grant_type;
  wire[3:0] T68;
  wire[3:0] T69;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[3:0] T80;
  wire T81;
  reg  init_sharer_cnt;
  wire T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[2:0] T89;
  wire T90;
  wire T91;
  wire[2:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg [25:0] xact_addr;
  wire[25:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[3:0] T105;
  wire[3:0] T106;
  wire[3:0] T107;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] T110;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T111;
  wire[5:0] T112;
  wire[5:0] T113;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T117;
  wire[511:0] T118;
  wire[511:0] T119;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T120;
  wire[3:0] T121;
  wire[3:0] T122;
  wire[3:0] T123;
  wire[3:0] outer_read_client_xact_id;
  wire[3:0] outer_write_rel_client_xact_id;
  wire[3:0] outer_write_acq_client_xact_id;
  wire[25:0] T124;
  wire[25:0] T125;
  wire[25:0] T126;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_write_acq_addr;
  wire T127;
  wire T128;
  wire T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[3:0] T145;
  wire[25:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  reg [1:0] probe_flags;
  wire[1:0] T150;
  wire[1:0] T151;
  wire[1:0] T152;
  wire[1:0] T153;
  wire[1:0] T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[3:0] T159;
  wire[3:0] T160;
  wire[3:0] T161;
  reg [3:0] xact_client_xact_id;
  wire[3:0] T162;
  wire[511:0] T163;
  wire[1:0] T164;
  reg  init_client_id;
  wire T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T100 & T1;
  assign T1 = state != 3'h0;
  assign T2 = reset ? 3'h0 : T3;
  assign T3 = T96 ? 3'h0 : T4;
  assign T4 = T94 ? T92 : T5;
  assign T5 = T90 ? T89 : T6;
  assign T6 = T87 ? T66 : T7;
  assign T7 = T64 ? T62 : T8;
  assign T8 = T32 ? T24 : T9;
  assign T9 = T22 ? T10 : state;
  assign T10 = T19 ? 3'h1 : T11;
  assign T11 = T14 ? 3'h3 : T12;
  assign T12 = T13 ? 3'h2 : 3'h4;
  assign T13 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T14 = T16 | T15;
  assign T15 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T16 = T18 | T17;
  assign T17 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T18 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T19 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T20;
  assign T20 = ~ T21;
  assign T21 = io_tile_incoherent | 2'h0;
  assign T22 = T23 & io_inner_acquire_valid;
  assign T23 = 3'h0 == state;
  assign T24 = pending_outer_write ? 3'h3 : T25;
  assign T25 = T26 ? 3'h2 : 3'h4;
  assign T26 = xact_a_type != 3'h3;
  assign T27 = T22 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T29 | T28;
  assign T28 = 3'h6 == xact_a_type;
  assign T29 = T31 | T30;
  assign T30 = 3'h5 == xact_a_type;
  assign T31 = 3'h3 == xact_a_type;
  assign T32 = T47 & T33;
  assign T33 = release_count == 1'h1;
  assign T34 = T35[1'h0:1'h0];
  assign T35 = reset ? 2'h0 : T36;
  assign T36 = T60 ? T58 : T37;
  assign T37 = T47 ? T45 : T38;
  assign T38 = T22 ? T40 : T39;
  assign T39 = {1'h0, release_count};
  assign T40 = T43 + T41;
  assign T41 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h1:1'h1];
  assign T43 = {1'h0, T44};
  assign T44 = probe_initial_flags[1'h0:1'h0];
  assign T45 = {1'h0, T46};
  assign T46 = release_count - 1'h1;
  assign T47 = T48 & io_outer_acquire_ready;
  assign T48 = T56 & T49;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T53 = T55 | T54;
  assign T54 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T55 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T56 = T57 & io_inner_release_valid;
  assign T57 = 3'h1 == state;
  assign T58 = {1'h0, T59};
  assign T59 = release_count - 1'h1;
  assign T60 = T56 & T61;
  assign T61 = T49 ^ 1'h1;
  assign T62 = pending_outer_write ? 3'h3 : T63;
  assign T63 = T26 ? 3'h2 : 3'h4;
  assign T64 = T60 & T65;
  assign T65 = release_count == 1'h1;
  assign T66 = T67 ? 3'h5 : 3'h0;
  assign T67 = grant_type != 4'h0;
  assign grant_type = T86 ? T80 : T68;
  assign T68 = T79 ? 4'h2 : T69;
  assign T69 = T78 ? 4'h3 : T70;
  assign T70 = T77 ? 4'h4 : T71;
  assign T71 = T76 ? 4'h6 : T72;
  assign T72 = T75 ? 4'h7 : T73;
  assign T73 = T74 ? 4'h8 : 4'h3;
  assign T74 = xact_a_type == 3'h6;
  assign T75 = xact_a_type == 3'h5;
  assign T76 = xact_a_type == 3'h4;
  assign T77 = xact_a_type == 3'h3;
  assign T78 = xact_a_type == 3'h2;
  assign T79 = xact_a_type == 3'h1;
  assign T80 = T81 ? 4'h1 : 4'h2;
  assign T81 = 1'h0 < init_sharer_cnt;
  assign T82 = T83[1'h0:1'h0];
  assign T83 = reset ? 2'h0 : T84;
  assign T84 = T22 ? 2'h2 : T85;
  assign T85 = {1'h0, init_sharer_cnt};
  assign T86 = xact_a_type == 3'h0;
  assign T87 = T88 & io_outer_acquire_ready;
  assign T88 = 3'h2 == state;
  assign T89 = T26 ? 3'h2 : 3'h4;
  assign T90 = T91 & io_outer_acquire_ready;
  assign T91 = 3'h3 == state;
  assign T92 = T93 ? 3'h5 : 3'h0;
  assign T93 = grant_type != 4'h0;
  assign T94 = T95 & io_inner_grant_ready;
  assign T95 = 3'h4 == state;
  assign T96 = T99 & T97;
  assign T97 = io_inner_finish_valid & T98;
  assign T98 = io_inner_finish_bits_payload_master_xact_id == 4'h1;
  assign T99 = 3'h5 == state;
  assign T100 = xact_addr == io_inner_release_bits_payload_addr;
  assign T101 = T22 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T102;
  assign T102 = T104 & T103;
  assign T103 = state != 3'h0;
  assign T104 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T105;
  assign T105 = T91 ? outer_write_acq_atomic_opcode : T106;
  assign T106 = T88 ? outer_read_atomic_opcode : T107;
  assign T107 = T48 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T108;
  assign T108 = T91 ? outer_write_acq_subword_addr : T109;
  assign T109 = T88 ? outer_read_subword_addr : T110;
  assign T110 = T48 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T111;
  assign T111 = T91 ? outer_write_acq_write_mask : T112;
  assign T112 = T88 ? outer_read_write_mask : T113;
  assign T113 = T48 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T114;
  assign T114 = T91 ? outer_write_acq_a_type : T115;
  assign T115 = T88 ? outer_read_a_type : T116;
  assign T116 = T48 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_read_a_type = 3'h2;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T117;
  assign T117 = T91 ? outer_write_acq_data : T118;
  assign T118 = T88 ? outer_read_data : T119;
  assign T119 = T48 ? outer_write_rel_data : outer_read_data;
  assign outer_read_data = 512'h0;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_write_acq_data = xact_data;
  assign T120 = T22 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T121;
  assign T121 = T91 ? outer_write_acq_client_xact_id : T122;
  assign T122 = T88 ? outer_read_client_xact_id : T123;
  assign T123 = T48 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_read_client_xact_id = 4'h1;
  assign outer_write_rel_client_xact_id = 4'h1;
  assign outer_write_acq_client_xact_id = 4'h1;
  assign io_outer_acquire_bits_payload_addr = T124;
  assign T124 = T91 ? outer_write_acq_addr : T125;
  assign T125 = T88 ? outer_read_addr : T126;
  assign T126 = T48 ? outer_write_rel_addr : outer_read_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T127;
  assign T127 = T91 ? 1'h1 : T128;
  assign T128 = T88 ? 1'h1 : T48;
  assign io_inner_release_ready = T129;
  assign T129 = T60 ? 1'h1 : T47;
  assign io_inner_probe_bits_payload_p_type = T130;
  assign T130 = T131;
  assign T131 = T144 ? 2'h1 : T132;
  assign T132 = T143 ? 2'h0 : T133;
  assign T133 = T142 ? 2'h2 : T134;
  assign T134 = T141 ? 2'h0 : T135;
  assign T135 = T140 ? 2'h2 : T136;
  assign T136 = T139 ? 2'h0 : T137;
  assign T137 = T138 ? 2'h0 : 2'h2;
  assign T138 = xact_a_type == 3'h6;
  assign T139 = xact_a_type == 3'h5;
  assign T140 = xact_a_type == 3'h4;
  assign T141 = xact_a_type == 3'h3;
  assign T142 = xact_a_type == 3'h2;
  assign T143 = xact_a_type == 3'h1;
  assign T144 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T145;
  assign T145 = 4'h1;
  assign io_inner_probe_bits_payload_addr = T146;
  assign T146 = xact_addr;
  assign io_inner_probe_bits_header_dst = T147;
  assign T147 = {1'h0, T148};
  assign T148 = T149 == 1'h0;
  assign T149 = probe_flags[1'h0:1'h0];
  assign T150 = reset ? 2'h0 : T151;
  assign T151 = T156 ? T153 : T152;
  assign T152 = T22 ? probe_initial_flags : probe_flags;
  assign T153 = probe_flags & T154;
  assign T154 = ~ T155;
  assign T155 = 1'h1 << T148;
  assign T156 = T57 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T157;
  assign T157 = T57 ? T158 : 1'h0;
  assign T158 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T159;
  assign T159 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T160;
  assign T160 = 4'h1;
  assign io_inner_grant_bits_payload_client_xact_id = T161;
  assign T161 = xact_client_xact_id;
  assign T162 = T22 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T163;
  assign T163 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T164;
  assign T164 = {1'h0, init_client_id};
  assign T165 = T166[1'h0:1'h0];
  assign T166 = reset ? 2'h0 : T167;
  assign T167 = T22 ? io_inner_acquire_bits_header_src : T168;
  assign T168 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T169;
  assign T169 = T170 ? 1'h1 : T95;
  assign T170 = T99 & T171;
  assign T171 = io_outer_grant_valid & T172;
  assign T172 = io_outer_grant_bits_payload_client_xact_id == 4'h1;
  assign io_inner_acquire_ready = T23;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T96) begin
      state <= 3'h0;
    end else if(T94) begin
      state <= T92;
    end else if(T90) begin
      state <= T89;
    end else if(T87) begin
      state <= T66;
    end else if(T64) begin
      state <= T62;
    end else if(T32) begin
      state <= T24;
    end else if(T22) begin
      state <= T10;
    end
    if(T22) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T34;
    init_sharer_cnt <= T82;
    if(T22) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T22) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T156) begin
      probe_flags <= T153;
    end else if(T22) begin
      probe_flags <= probe_initial_flags;
    end
    if(T22) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T165;
  end
endmodule

module AcquireTracker_1(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [3:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[3:0] io_inner_grant_bits_payload_client_xact_id,
    output[3:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [3:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[3:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [3:0] io_inner_release_bits_payload_client_xact_id,
    input [3:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[3:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [3:0] io_outer_grant_bits_payload_client_xact_id,
    input [3:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[3:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] probe_initial_flags;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  reg [2:0] xact_a_type;
  wire[2:0] T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  reg  release_count;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[2:0] T62;
  wire[2:0] T63;
  wire T64;
  wire T65;
  wire[2:0] T66;
  wire T67;
  wire[3:0] grant_type;
  wire[3:0] T68;
  wire[3:0] T69;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[3:0] T80;
  wire T81;
  reg  init_sharer_cnt;
  wire T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[2:0] T89;
  wire T90;
  wire T91;
  wire[2:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg [25:0] xact_addr;
  wire[25:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[3:0] T105;
  wire[3:0] T106;
  wire[3:0] T107;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] T110;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T111;
  wire[5:0] T112;
  wire[5:0] T113;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T117;
  wire[511:0] T118;
  wire[511:0] T119;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T120;
  wire[3:0] T121;
  wire[3:0] T122;
  wire[3:0] T123;
  wire[3:0] outer_read_client_xact_id;
  wire[3:0] outer_write_rel_client_xact_id;
  wire[3:0] outer_write_acq_client_xact_id;
  wire[25:0] T124;
  wire[25:0] T125;
  wire[25:0] T126;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_write_acq_addr;
  wire T127;
  wire T128;
  wire T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[3:0] T145;
  wire[25:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  reg [1:0] probe_flags;
  wire[1:0] T150;
  wire[1:0] T151;
  wire[1:0] T152;
  wire[1:0] T153;
  wire[1:0] T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[3:0] T159;
  wire[3:0] T160;
  wire[3:0] T161;
  reg [3:0] xact_client_xact_id;
  wire[3:0] T162;
  wire[511:0] T163;
  wire[1:0] T164;
  reg  init_client_id;
  wire T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T100 & T1;
  assign T1 = state != 3'h0;
  assign T2 = reset ? 3'h0 : T3;
  assign T3 = T96 ? 3'h0 : T4;
  assign T4 = T94 ? T92 : T5;
  assign T5 = T90 ? T89 : T6;
  assign T6 = T87 ? T66 : T7;
  assign T7 = T64 ? T62 : T8;
  assign T8 = T32 ? T24 : T9;
  assign T9 = T22 ? T10 : state;
  assign T10 = T19 ? 3'h1 : T11;
  assign T11 = T14 ? 3'h3 : T12;
  assign T12 = T13 ? 3'h2 : 3'h4;
  assign T13 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T14 = T16 | T15;
  assign T15 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T16 = T18 | T17;
  assign T17 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T18 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T19 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T20;
  assign T20 = ~ T21;
  assign T21 = io_tile_incoherent | 2'h0;
  assign T22 = T23 & io_inner_acquire_valid;
  assign T23 = 3'h0 == state;
  assign T24 = pending_outer_write ? 3'h3 : T25;
  assign T25 = T26 ? 3'h2 : 3'h4;
  assign T26 = xact_a_type != 3'h3;
  assign T27 = T22 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T29 | T28;
  assign T28 = 3'h6 == xact_a_type;
  assign T29 = T31 | T30;
  assign T30 = 3'h5 == xact_a_type;
  assign T31 = 3'h3 == xact_a_type;
  assign T32 = T47 & T33;
  assign T33 = release_count == 1'h1;
  assign T34 = T35[1'h0:1'h0];
  assign T35 = reset ? 2'h0 : T36;
  assign T36 = T60 ? T58 : T37;
  assign T37 = T47 ? T45 : T38;
  assign T38 = T22 ? T40 : T39;
  assign T39 = {1'h0, release_count};
  assign T40 = T43 + T41;
  assign T41 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h1:1'h1];
  assign T43 = {1'h0, T44};
  assign T44 = probe_initial_flags[1'h0:1'h0];
  assign T45 = {1'h0, T46};
  assign T46 = release_count - 1'h1;
  assign T47 = T48 & io_outer_acquire_ready;
  assign T48 = T56 & T49;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T53 = T55 | T54;
  assign T54 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T55 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T56 = T57 & io_inner_release_valid;
  assign T57 = 3'h1 == state;
  assign T58 = {1'h0, T59};
  assign T59 = release_count - 1'h1;
  assign T60 = T56 & T61;
  assign T61 = T49 ^ 1'h1;
  assign T62 = pending_outer_write ? 3'h3 : T63;
  assign T63 = T26 ? 3'h2 : 3'h4;
  assign T64 = T60 & T65;
  assign T65 = release_count == 1'h1;
  assign T66 = T67 ? 3'h5 : 3'h0;
  assign T67 = grant_type != 4'h0;
  assign grant_type = T86 ? T80 : T68;
  assign T68 = T79 ? 4'h2 : T69;
  assign T69 = T78 ? 4'h3 : T70;
  assign T70 = T77 ? 4'h4 : T71;
  assign T71 = T76 ? 4'h6 : T72;
  assign T72 = T75 ? 4'h7 : T73;
  assign T73 = T74 ? 4'h8 : 4'h3;
  assign T74 = xact_a_type == 3'h6;
  assign T75 = xact_a_type == 3'h5;
  assign T76 = xact_a_type == 3'h4;
  assign T77 = xact_a_type == 3'h3;
  assign T78 = xact_a_type == 3'h2;
  assign T79 = xact_a_type == 3'h1;
  assign T80 = T81 ? 4'h1 : 4'h2;
  assign T81 = 1'h0 < init_sharer_cnt;
  assign T82 = T83[1'h0:1'h0];
  assign T83 = reset ? 2'h0 : T84;
  assign T84 = T22 ? 2'h2 : T85;
  assign T85 = {1'h0, init_sharer_cnt};
  assign T86 = xact_a_type == 3'h0;
  assign T87 = T88 & io_outer_acquire_ready;
  assign T88 = 3'h2 == state;
  assign T89 = T26 ? 3'h2 : 3'h4;
  assign T90 = T91 & io_outer_acquire_ready;
  assign T91 = 3'h3 == state;
  assign T92 = T93 ? 3'h5 : 3'h0;
  assign T93 = grant_type != 4'h0;
  assign T94 = T95 & io_inner_grant_ready;
  assign T95 = 3'h4 == state;
  assign T96 = T99 & T97;
  assign T97 = io_inner_finish_valid & T98;
  assign T98 = io_inner_finish_bits_payload_master_xact_id == 4'h2;
  assign T99 = 3'h5 == state;
  assign T100 = xact_addr == io_inner_release_bits_payload_addr;
  assign T101 = T22 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T102;
  assign T102 = T104 & T103;
  assign T103 = state != 3'h0;
  assign T104 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T105;
  assign T105 = T91 ? outer_write_acq_atomic_opcode : T106;
  assign T106 = T88 ? outer_read_atomic_opcode : T107;
  assign T107 = T48 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T108;
  assign T108 = T91 ? outer_write_acq_subword_addr : T109;
  assign T109 = T88 ? outer_read_subword_addr : T110;
  assign T110 = T48 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T111;
  assign T111 = T91 ? outer_write_acq_write_mask : T112;
  assign T112 = T88 ? outer_read_write_mask : T113;
  assign T113 = T48 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T114;
  assign T114 = T91 ? outer_write_acq_a_type : T115;
  assign T115 = T88 ? outer_read_a_type : T116;
  assign T116 = T48 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_read_a_type = 3'h2;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T117;
  assign T117 = T91 ? outer_write_acq_data : T118;
  assign T118 = T88 ? outer_read_data : T119;
  assign T119 = T48 ? outer_write_rel_data : outer_read_data;
  assign outer_read_data = 512'h0;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_write_acq_data = xact_data;
  assign T120 = T22 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T121;
  assign T121 = T91 ? outer_write_acq_client_xact_id : T122;
  assign T122 = T88 ? outer_read_client_xact_id : T123;
  assign T123 = T48 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_read_client_xact_id = 4'h2;
  assign outer_write_rel_client_xact_id = 4'h2;
  assign outer_write_acq_client_xact_id = 4'h2;
  assign io_outer_acquire_bits_payload_addr = T124;
  assign T124 = T91 ? outer_write_acq_addr : T125;
  assign T125 = T88 ? outer_read_addr : T126;
  assign T126 = T48 ? outer_write_rel_addr : outer_read_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T127;
  assign T127 = T91 ? 1'h1 : T128;
  assign T128 = T88 ? 1'h1 : T48;
  assign io_inner_release_ready = T129;
  assign T129 = T60 ? 1'h1 : T47;
  assign io_inner_probe_bits_payload_p_type = T130;
  assign T130 = T131;
  assign T131 = T144 ? 2'h1 : T132;
  assign T132 = T143 ? 2'h0 : T133;
  assign T133 = T142 ? 2'h2 : T134;
  assign T134 = T141 ? 2'h0 : T135;
  assign T135 = T140 ? 2'h2 : T136;
  assign T136 = T139 ? 2'h0 : T137;
  assign T137 = T138 ? 2'h0 : 2'h2;
  assign T138 = xact_a_type == 3'h6;
  assign T139 = xact_a_type == 3'h5;
  assign T140 = xact_a_type == 3'h4;
  assign T141 = xact_a_type == 3'h3;
  assign T142 = xact_a_type == 3'h2;
  assign T143 = xact_a_type == 3'h1;
  assign T144 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T145;
  assign T145 = 4'h2;
  assign io_inner_probe_bits_payload_addr = T146;
  assign T146 = xact_addr;
  assign io_inner_probe_bits_header_dst = T147;
  assign T147 = {1'h0, T148};
  assign T148 = T149 == 1'h0;
  assign T149 = probe_flags[1'h0:1'h0];
  assign T150 = reset ? 2'h0 : T151;
  assign T151 = T156 ? T153 : T152;
  assign T152 = T22 ? probe_initial_flags : probe_flags;
  assign T153 = probe_flags & T154;
  assign T154 = ~ T155;
  assign T155 = 1'h1 << T148;
  assign T156 = T57 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T157;
  assign T157 = T57 ? T158 : 1'h0;
  assign T158 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T159;
  assign T159 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T160;
  assign T160 = 4'h2;
  assign io_inner_grant_bits_payload_client_xact_id = T161;
  assign T161 = xact_client_xact_id;
  assign T162 = T22 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T163;
  assign T163 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T164;
  assign T164 = {1'h0, init_client_id};
  assign T165 = T166[1'h0:1'h0];
  assign T166 = reset ? 2'h0 : T167;
  assign T167 = T22 ? io_inner_acquire_bits_header_src : T168;
  assign T168 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T169;
  assign T169 = T170 ? 1'h1 : T95;
  assign T170 = T99 & T171;
  assign T171 = io_outer_grant_valid & T172;
  assign T172 = io_outer_grant_bits_payload_client_xact_id == 4'h2;
  assign io_inner_acquire_ready = T23;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T96) begin
      state <= 3'h0;
    end else if(T94) begin
      state <= T92;
    end else if(T90) begin
      state <= T89;
    end else if(T87) begin
      state <= T66;
    end else if(T64) begin
      state <= T62;
    end else if(T32) begin
      state <= T24;
    end else if(T22) begin
      state <= T10;
    end
    if(T22) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T34;
    init_sharer_cnt <= T82;
    if(T22) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T22) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T156) begin
      probe_flags <= T153;
    end else if(T22) begin
      probe_flags <= probe_initial_flags;
    end
    if(T22) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T165;
  end
endmodule

module AcquireTracker_2(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [3:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[3:0] io_inner_grant_bits_payload_client_xact_id,
    output[3:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [3:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[3:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [3:0] io_inner_release_bits_payload_client_xact_id,
    input [3:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[3:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [3:0] io_outer_grant_bits_payload_client_xact_id,
    input [3:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[3:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] probe_initial_flags;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  reg [2:0] xact_a_type;
  wire[2:0] T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  reg  release_count;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[2:0] T62;
  wire[2:0] T63;
  wire T64;
  wire T65;
  wire[2:0] T66;
  wire T67;
  wire[3:0] grant_type;
  wire[3:0] T68;
  wire[3:0] T69;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[3:0] T80;
  wire T81;
  reg  init_sharer_cnt;
  wire T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[2:0] T89;
  wire T90;
  wire T91;
  wire[2:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg [25:0] xact_addr;
  wire[25:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[3:0] T105;
  wire[3:0] T106;
  wire[3:0] T107;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] T110;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T111;
  wire[5:0] T112;
  wire[5:0] T113;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T117;
  wire[511:0] T118;
  wire[511:0] T119;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T120;
  wire[3:0] T121;
  wire[3:0] T122;
  wire[3:0] T123;
  wire[3:0] outer_read_client_xact_id;
  wire[3:0] outer_write_rel_client_xact_id;
  wire[3:0] outer_write_acq_client_xact_id;
  wire[25:0] T124;
  wire[25:0] T125;
  wire[25:0] T126;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_write_acq_addr;
  wire T127;
  wire T128;
  wire T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[3:0] T145;
  wire[25:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  reg [1:0] probe_flags;
  wire[1:0] T150;
  wire[1:0] T151;
  wire[1:0] T152;
  wire[1:0] T153;
  wire[1:0] T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[3:0] T159;
  wire[3:0] T160;
  wire[3:0] T161;
  reg [3:0] xact_client_xact_id;
  wire[3:0] T162;
  wire[511:0] T163;
  wire[1:0] T164;
  reg  init_client_id;
  wire T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T100 & T1;
  assign T1 = state != 3'h0;
  assign T2 = reset ? 3'h0 : T3;
  assign T3 = T96 ? 3'h0 : T4;
  assign T4 = T94 ? T92 : T5;
  assign T5 = T90 ? T89 : T6;
  assign T6 = T87 ? T66 : T7;
  assign T7 = T64 ? T62 : T8;
  assign T8 = T32 ? T24 : T9;
  assign T9 = T22 ? T10 : state;
  assign T10 = T19 ? 3'h1 : T11;
  assign T11 = T14 ? 3'h3 : T12;
  assign T12 = T13 ? 3'h2 : 3'h4;
  assign T13 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T14 = T16 | T15;
  assign T15 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T16 = T18 | T17;
  assign T17 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T18 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T19 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T20;
  assign T20 = ~ T21;
  assign T21 = io_tile_incoherent | 2'h0;
  assign T22 = T23 & io_inner_acquire_valid;
  assign T23 = 3'h0 == state;
  assign T24 = pending_outer_write ? 3'h3 : T25;
  assign T25 = T26 ? 3'h2 : 3'h4;
  assign T26 = xact_a_type != 3'h3;
  assign T27 = T22 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T29 | T28;
  assign T28 = 3'h6 == xact_a_type;
  assign T29 = T31 | T30;
  assign T30 = 3'h5 == xact_a_type;
  assign T31 = 3'h3 == xact_a_type;
  assign T32 = T47 & T33;
  assign T33 = release_count == 1'h1;
  assign T34 = T35[1'h0:1'h0];
  assign T35 = reset ? 2'h0 : T36;
  assign T36 = T60 ? T58 : T37;
  assign T37 = T47 ? T45 : T38;
  assign T38 = T22 ? T40 : T39;
  assign T39 = {1'h0, release_count};
  assign T40 = T43 + T41;
  assign T41 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h1:1'h1];
  assign T43 = {1'h0, T44};
  assign T44 = probe_initial_flags[1'h0:1'h0];
  assign T45 = {1'h0, T46};
  assign T46 = release_count - 1'h1;
  assign T47 = T48 & io_outer_acquire_ready;
  assign T48 = T56 & T49;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T53 = T55 | T54;
  assign T54 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T55 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T56 = T57 & io_inner_release_valid;
  assign T57 = 3'h1 == state;
  assign T58 = {1'h0, T59};
  assign T59 = release_count - 1'h1;
  assign T60 = T56 & T61;
  assign T61 = T49 ^ 1'h1;
  assign T62 = pending_outer_write ? 3'h3 : T63;
  assign T63 = T26 ? 3'h2 : 3'h4;
  assign T64 = T60 & T65;
  assign T65 = release_count == 1'h1;
  assign T66 = T67 ? 3'h5 : 3'h0;
  assign T67 = grant_type != 4'h0;
  assign grant_type = T86 ? T80 : T68;
  assign T68 = T79 ? 4'h2 : T69;
  assign T69 = T78 ? 4'h3 : T70;
  assign T70 = T77 ? 4'h4 : T71;
  assign T71 = T76 ? 4'h6 : T72;
  assign T72 = T75 ? 4'h7 : T73;
  assign T73 = T74 ? 4'h8 : 4'h3;
  assign T74 = xact_a_type == 3'h6;
  assign T75 = xact_a_type == 3'h5;
  assign T76 = xact_a_type == 3'h4;
  assign T77 = xact_a_type == 3'h3;
  assign T78 = xact_a_type == 3'h2;
  assign T79 = xact_a_type == 3'h1;
  assign T80 = T81 ? 4'h1 : 4'h2;
  assign T81 = 1'h0 < init_sharer_cnt;
  assign T82 = T83[1'h0:1'h0];
  assign T83 = reset ? 2'h0 : T84;
  assign T84 = T22 ? 2'h2 : T85;
  assign T85 = {1'h0, init_sharer_cnt};
  assign T86 = xact_a_type == 3'h0;
  assign T87 = T88 & io_outer_acquire_ready;
  assign T88 = 3'h2 == state;
  assign T89 = T26 ? 3'h2 : 3'h4;
  assign T90 = T91 & io_outer_acquire_ready;
  assign T91 = 3'h3 == state;
  assign T92 = T93 ? 3'h5 : 3'h0;
  assign T93 = grant_type != 4'h0;
  assign T94 = T95 & io_inner_grant_ready;
  assign T95 = 3'h4 == state;
  assign T96 = T99 & T97;
  assign T97 = io_inner_finish_valid & T98;
  assign T98 = io_inner_finish_bits_payload_master_xact_id == 4'h3;
  assign T99 = 3'h5 == state;
  assign T100 = xact_addr == io_inner_release_bits_payload_addr;
  assign T101 = T22 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T102;
  assign T102 = T104 & T103;
  assign T103 = state != 3'h0;
  assign T104 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T105;
  assign T105 = T91 ? outer_write_acq_atomic_opcode : T106;
  assign T106 = T88 ? outer_read_atomic_opcode : T107;
  assign T107 = T48 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T108;
  assign T108 = T91 ? outer_write_acq_subword_addr : T109;
  assign T109 = T88 ? outer_read_subword_addr : T110;
  assign T110 = T48 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T111;
  assign T111 = T91 ? outer_write_acq_write_mask : T112;
  assign T112 = T88 ? outer_read_write_mask : T113;
  assign T113 = T48 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T114;
  assign T114 = T91 ? outer_write_acq_a_type : T115;
  assign T115 = T88 ? outer_read_a_type : T116;
  assign T116 = T48 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_read_a_type = 3'h2;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T117;
  assign T117 = T91 ? outer_write_acq_data : T118;
  assign T118 = T88 ? outer_read_data : T119;
  assign T119 = T48 ? outer_write_rel_data : outer_read_data;
  assign outer_read_data = 512'h0;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_write_acq_data = xact_data;
  assign T120 = T22 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T121;
  assign T121 = T91 ? outer_write_acq_client_xact_id : T122;
  assign T122 = T88 ? outer_read_client_xact_id : T123;
  assign T123 = T48 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_read_client_xact_id = 4'h3;
  assign outer_write_rel_client_xact_id = 4'h3;
  assign outer_write_acq_client_xact_id = 4'h3;
  assign io_outer_acquire_bits_payload_addr = T124;
  assign T124 = T91 ? outer_write_acq_addr : T125;
  assign T125 = T88 ? outer_read_addr : T126;
  assign T126 = T48 ? outer_write_rel_addr : outer_read_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T127;
  assign T127 = T91 ? 1'h1 : T128;
  assign T128 = T88 ? 1'h1 : T48;
  assign io_inner_release_ready = T129;
  assign T129 = T60 ? 1'h1 : T47;
  assign io_inner_probe_bits_payload_p_type = T130;
  assign T130 = T131;
  assign T131 = T144 ? 2'h1 : T132;
  assign T132 = T143 ? 2'h0 : T133;
  assign T133 = T142 ? 2'h2 : T134;
  assign T134 = T141 ? 2'h0 : T135;
  assign T135 = T140 ? 2'h2 : T136;
  assign T136 = T139 ? 2'h0 : T137;
  assign T137 = T138 ? 2'h0 : 2'h2;
  assign T138 = xact_a_type == 3'h6;
  assign T139 = xact_a_type == 3'h5;
  assign T140 = xact_a_type == 3'h4;
  assign T141 = xact_a_type == 3'h3;
  assign T142 = xact_a_type == 3'h2;
  assign T143 = xact_a_type == 3'h1;
  assign T144 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T145;
  assign T145 = 4'h3;
  assign io_inner_probe_bits_payload_addr = T146;
  assign T146 = xact_addr;
  assign io_inner_probe_bits_header_dst = T147;
  assign T147 = {1'h0, T148};
  assign T148 = T149 == 1'h0;
  assign T149 = probe_flags[1'h0:1'h0];
  assign T150 = reset ? 2'h0 : T151;
  assign T151 = T156 ? T153 : T152;
  assign T152 = T22 ? probe_initial_flags : probe_flags;
  assign T153 = probe_flags & T154;
  assign T154 = ~ T155;
  assign T155 = 1'h1 << T148;
  assign T156 = T57 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T157;
  assign T157 = T57 ? T158 : 1'h0;
  assign T158 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T159;
  assign T159 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T160;
  assign T160 = 4'h3;
  assign io_inner_grant_bits_payload_client_xact_id = T161;
  assign T161 = xact_client_xact_id;
  assign T162 = T22 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T163;
  assign T163 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T164;
  assign T164 = {1'h0, init_client_id};
  assign T165 = T166[1'h0:1'h0];
  assign T166 = reset ? 2'h0 : T167;
  assign T167 = T22 ? io_inner_acquire_bits_header_src : T168;
  assign T168 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T169;
  assign T169 = T170 ? 1'h1 : T95;
  assign T170 = T99 & T171;
  assign T171 = io_outer_grant_valid & T172;
  assign T172 = io_outer_grant_bits_payload_client_xact_id == 4'h3;
  assign io_inner_acquire_ready = T23;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T96) begin
      state <= 3'h0;
    end else if(T94) begin
      state <= T92;
    end else if(T90) begin
      state <= T89;
    end else if(T87) begin
      state <= T66;
    end else if(T64) begin
      state <= T62;
    end else if(T32) begin
      state <= T24;
    end else if(T22) begin
      state <= T10;
    end
    if(T22) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T34;
    init_sharer_cnt <= T82;
    if(T22) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T22) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T156) begin
      probe_flags <= T153;
    end else if(T22) begin
      probe_flags <= probe_initial_flags;
    end
    if(T22) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T165;
  end
endmodule

module AcquireTracker_3(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [3:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[3:0] io_inner_grant_bits_payload_client_xact_id,
    output[3:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [3:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[3:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [3:0] io_inner_release_bits_payload_client_xact_id,
    input [3:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[3:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [3:0] io_outer_grant_bits_payload_client_xact_id,
    input [3:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[3:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] probe_initial_flags;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  reg [2:0] xact_a_type;
  wire[2:0] T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  reg  release_count;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[2:0] T62;
  wire[2:0] T63;
  wire T64;
  wire T65;
  wire[2:0] T66;
  wire T67;
  wire[3:0] grant_type;
  wire[3:0] T68;
  wire[3:0] T69;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[3:0] T80;
  wire T81;
  reg  init_sharer_cnt;
  wire T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[2:0] T89;
  wire T90;
  wire T91;
  wire[2:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg [25:0] xact_addr;
  wire[25:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[3:0] T105;
  wire[3:0] T106;
  wire[3:0] T107;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] T110;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T111;
  wire[5:0] T112;
  wire[5:0] T113;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T117;
  wire[511:0] T118;
  wire[511:0] T119;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T120;
  wire[3:0] T121;
  wire[3:0] T122;
  wire[3:0] T123;
  wire[3:0] outer_read_client_xact_id;
  wire[3:0] outer_write_rel_client_xact_id;
  wire[3:0] outer_write_acq_client_xact_id;
  wire[25:0] T124;
  wire[25:0] T125;
  wire[25:0] T126;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_write_acq_addr;
  wire T127;
  wire T128;
  wire T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[3:0] T145;
  wire[25:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  reg [1:0] probe_flags;
  wire[1:0] T150;
  wire[1:0] T151;
  wire[1:0] T152;
  wire[1:0] T153;
  wire[1:0] T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[3:0] T159;
  wire[3:0] T160;
  wire[3:0] T161;
  reg [3:0] xact_client_xact_id;
  wire[3:0] T162;
  wire[511:0] T163;
  wire[1:0] T164;
  reg  init_client_id;
  wire T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T100 & T1;
  assign T1 = state != 3'h0;
  assign T2 = reset ? 3'h0 : T3;
  assign T3 = T96 ? 3'h0 : T4;
  assign T4 = T94 ? T92 : T5;
  assign T5 = T90 ? T89 : T6;
  assign T6 = T87 ? T66 : T7;
  assign T7 = T64 ? T62 : T8;
  assign T8 = T32 ? T24 : T9;
  assign T9 = T22 ? T10 : state;
  assign T10 = T19 ? 3'h1 : T11;
  assign T11 = T14 ? 3'h3 : T12;
  assign T12 = T13 ? 3'h2 : 3'h4;
  assign T13 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T14 = T16 | T15;
  assign T15 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T16 = T18 | T17;
  assign T17 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T18 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T19 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T20;
  assign T20 = ~ T21;
  assign T21 = io_tile_incoherent | 2'h0;
  assign T22 = T23 & io_inner_acquire_valid;
  assign T23 = 3'h0 == state;
  assign T24 = pending_outer_write ? 3'h3 : T25;
  assign T25 = T26 ? 3'h2 : 3'h4;
  assign T26 = xact_a_type != 3'h3;
  assign T27 = T22 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T29 | T28;
  assign T28 = 3'h6 == xact_a_type;
  assign T29 = T31 | T30;
  assign T30 = 3'h5 == xact_a_type;
  assign T31 = 3'h3 == xact_a_type;
  assign T32 = T47 & T33;
  assign T33 = release_count == 1'h1;
  assign T34 = T35[1'h0:1'h0];
  assign T35 = reset ? 2'h0 : T36;
  assign T36 = T60 ? T58 : T37;
  assign T37 = T47 ? T45 : T38;
  assign T38 = T22 ? T40 : T39;
  assign T39 = {1'h0, release_count};
  assign T40 = T43 + T41;
  assign T41 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h1:1'h1];
  assign T43 = {1'h0, T44};
  assign T44 = probe_initial_flags[1'h0:1'h0];
  assign T45 = {1'h0, T46};
  assign T46 = release_count - 1'h1;
  assign T47 = T48 & io_outer_acquire_ready;
  assign T48 = T56 & T49;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T53 = T55 | T54;
  assign T54 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T55 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T56 = T57 & io_inner_release_valid;
  assign T57 = 3'h1 == state;
  assign T58 = {1'h0, T59};
  assign T59 = release_count - 1'h1;
  assign T60 = T56 & T61;
  assign T61 = T49 ^ 1'h1;
  assign T62 = pending_outer_write ? 3'h3 : T63;
  assign T63 = T26 ? 3'h2 : 3'h4;
  assign T64 = T60 & T65;
  assign T65 = release_count == 1'h1;
  assign T66 = T67 ? 3'h5 : 3'h0;
  assign T67 = grant_type != 4'h0;
  assign grant_type = T86 ? T80 : T68;
  assign T68 = T79 ? 4'h2 : T69;
  assign T69 = T78 ? 4'h3 : T70;
  assign T70 = T77 ? 4'h4 : T71;
  assign T71 = T76 ? 4'h6 : T72;
  assign T72 = T75 ? 4'h7 : T73;
  assign T73 = T74 ? 4'h8 : 4'h3;
  assign T74 = xact_a_type == 3'h6;
  assign T75 = xact_a_type == 3'h5;
  assign T76 = xact_a_type == 3'h4;
  assign T77 = xact_a_type == 3'h3;
  assign T78 = xact_a_type == 3'h2;
  assign T79 = xact_a_type == 3'h1;
  assign T80 = T81 ? 4'h1 : 4'h2;
  assign T81 = 1'h0 < init_sharer_cnt;
  assign T82 = T83[1'h0:1'h0];
  assign T83 = reset ? 2'h0 : T84;
  assign T84 = T22 ? 2'h2 : T85;
  assign T85 = {1'h0, init_sharer_cnt};
  assign T86 = xact_a_type == 3'h0;
  assign T87 = T88 & io_outer_acquire_ready;
  assign T88 = 3'h2 == state;
  assign T89 = T26 ? 3'h2 : 3'h4;
  assign T90 = T91 & io_outer_acquire_ready;
  assign T91 = 3'h3 == state;
  assign T92 = T93 ? 3'h5 : 3'h0;
  assign T93 = grant_type != 4'h0;
  assign T94 = T95 & io_inner_grant_ready;
  assign T95 = 3'h4 == state;
  assign T96 = T99 & T97;
  assign T97 = io_inner_finish_valid & T98;
  assign T98 = io_inner_finish_bits_payload_master_xact_id == 4'h4;
  assign T99 = 3'h5 == state;
  assign T100 = xact_addr == io_inner_release_bits_payload_addr;
  assign T101 = T22 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T102;
  assign T102 = T104 & T103;
  assign T103 = state != 3'h0;
  assign T104 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T105;
  assign T105 = T91 ? outer_write_acq_atomic_opcode : T106;
  assign T106 = T88 ? outer_read_atomic_opcode : T107;
  assign T107 = T48 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T108;
  assign T108 = T91 ? outer_write_acq_subword_addr : T109;
  assign T109 = T88 ? outer_read_subword_addr : T110;
  assign T110 = T48 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T111;
  assign T111 = T91 ? outer_write_acq_write_mask : T112;
  assign T112 = T88 ? outer_read_write_mask : T113;
  assign T113 = T48 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T114;
  assign T114 = T91 ? outer_write_acq_a_type : T115;
  assign T115 = T88 ? outer_read_a_type : T116;
  assign T116 = T48 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_read_a_type = 3'h2;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T117;
  assign T117 = T91 ? outer_write_acq_data : T118;
  assign T118 = T88 ? outer_read_data : T119;
  assign T119 = T48 ? outer_write_rel_data : outer_read_data;
  assign outer_read_data = 512'h0;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_write_acq_data = xact_data;
  assign T120 = T22 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T121;
  assign T121 = T91 ? outer_write_acq_client_xact_id : T122;
  assign T122 = T88 ? outer_read_client_xact_id : T123;
  assign T123 = T48 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_read_client_xact_id = 4'h4;
  assign outer_write_rel_client_xact_id = 4'h4;
  assign outer_write_acq_client_xact_id = 4'h4;
  assign io_outer_acquire_bits_payload_addr = T124;
  assign T124 = T91 ? outer_write_acq_addr : T125;
  assign T125 = T88 ? outer_read_addr : T126;
  assign T126 = T48 ? outer_write_rel_addr : outer_read_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T127;
  assign T127 = T91 ? 1'h1 : T128;
  assign T128 = T88 ? 1'h1 : T48;
  assign io_inner_release_ready = T129;
  assign T129 = T60 ? 1'h1 : T47;
  assign io_inner_probe_bits_payload_p_type = T130;
  assign T130 = T131;
  assign T131 = T144 ? 2'h1 : T132;
  assign T132 = T143 ? 2'h0 : T133;
  assign T133 = T142 ? 2'h2 : T134;
  assign T134 = T141 ? 2'h0 : T135;
  assign T135 = T140 ? 2'h2 : T136;
  assign T136 = T139 ? 2'h0 : T137;
  assign T137 = T138 ? 2'h0 : 2'h2;
  assign T138 = xact_a_type == 3'h6;
  assign T139 = xact_a_type == 3'h5;
  assign T140 = xact_a_type == 3'h4;
  assign T141 = xact_a_type == 3'h3;
  assign T142 = xact_a_type == 3'h2;
  assign T143 = xact_a_type == 3'h1;
  assign T144 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T145;
  assign T145 = 4'h4;
  assign io_inner_probe_bits_payload_addr = T146;
  assign T146 = xact_addr;
  assign io_inner_probe_bits_header_dst = T147;
  assign T147 = {1'h0, T148};
  assign T148 = T149 == 1'h0;
  assign T149 = probe_flags[1'h0:1'h0];
  assign T150 = reset ? 2'h0 : T151;
  assign T151 = T156 ? T153 : T152;
  assign T152 = T22 ? probe_initial_flags : probe_flags;
  assign T153 = probe_flags & T154;
  assign T154 = ~ T155;
  assign T155 = 1'h1 << T148;
  assign T156 = T57 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T157;
  assign T157 = T57 ? T158 : 1'h0;
  assign T158 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T159;
  assign T159 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T160;
  assign T160 = 4'h4;
  assign io_inner_grant_bits_payload_client_xact_id = T161;
  assign T161 = xact_client_xact_id;
  assign T162 = T22 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T163;
  assign T163 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T164;
  assign T164 = {1'h0, init_client_id};
  assign T165 = T166[1'h0:1'h0];
  assign T166 = reset ? 2'h0 : T167;
  assign T167 = T22 ? io_inner_acquire_bits_header_src : T168;
  assign T168 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T169;
  assign T169 = T170 ? 1'h1 : T95;
  assign T170 = T99 & T171;
  assign T171 = io_outer_grant_valid & T172;
  assign T172 = io_outer_grant_bits_payload_client_xact_id == 4'h4;
  assign io_inner_acquire_ready = T23;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T96) begin
      state <= 3'h0;
    end else if(T94) begin
      state <= T92;
    end else if(T90) begin
      state <= T89;
    end else if(T87) begin
      state <= T66;
    end else if(T64) begin
      state <= T62;
    end else if(T32) begin
      state <= T24;
    end else if(T22) begin
      state <= T10;
    end
    if(T22) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T34;
    init_sharer_cnt <= T82;
    if(T22) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T22) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T156) begin
      probe_flags <= T153;
    end else if(T22) begin
      probe_flags <= probe_initial_flags;
    end
    if(T22) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T165;
  end
endmodule

module Arbiter_11(
    output io_in_4_ready,
    input  io_in_4_valid,
    input  io_in_4_bits,
    output io_in_3_ready,
    input  io_in_3_valid,
    input  io_in_3_bits,
    output io_in_2_ready,
    input  io_in_2_valid,
    input  io_in_2_bits,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire[2:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : 3'h4;
  assign io_out_bits = T5;
  assign T5 = T13 ? io_in_4_bits : T6;
  assign T6 = T12 ? T10 : T7;
  assign T7 = T8 ? io_in_1_bits : io_in_0_bits;
  assign T8 = T9[1'h0:1'h0];
  assign T9 = T0;
  assign T10 = T11 ? io_in_3_bits : io_in_2_bits;
  assign T11 = T9[1'h0:1'h0];
  assign T12 = T9[1'h1:1'h1];
  assign T13 = T9[2'h2:2'h2];
  assign io_out_valid = T14;
  assign T14 = T21 ? io_in_4_valid : T15;
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? io_in_1_valid : io_in_0_valid;
  assign T17 = T9[1'h0:1'h0];
  assign T18 = T19 ? io_in_3_valid : io_in_2_valid;
  assign T19 = T9[1'h0:1'h0];
  assign T20 = T9[1'h1:1'h1];
  assign T21 = T9[2'h2:2'h2];
  assign io_in_0_ready = T22;
  assign T22 = T23 & io_out_ready;
  assign T23 = 1'h1;
  assign io_in_1_ready = T24;
  assign T24 = T25 & io_out_ready;
  assign T25 = T26;
  assign T26 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T27;
  assign T27 = T28 & io_out_ready;
  assign T28 = T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T31;
  assign T31 = T32 & io_out_ready;
  assign T32 = T33;
  assign T33 = T34 ^ 1'h1;
  assign T34 = T35 | io_in_2_valid;
  assign T35 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T36;
  assign T36 = T37 & io_out_ready;
  assign T37 = T38;
  assign T38 = T39 ^ 1'h1;
  assign T39 = T40 | io_in_3_valid;
  assign T40 = T41 | io_in_2_valid;
  assign T41 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_12(
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr,
    input [3:0] io_in_4_bits_payload_master_xact_id,
    input [1:0] io_in_4_bits_payload_p_type,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr,
    input [3:0] io_in_3_bits_payload_master_xact_id,
    input [1:0] io_in_3_bits_payload_p_type,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [3:0] io_in_2_bits_payload_master_xact_id,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [3:0] io_in_1_bits_payload_master_xact_id,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [3:0] io_in_0_bits_payload_master_xact_id,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[3:0] io_out_bits_payload_master_xact_id,
    output[1:0] io_out_bits_payload_p_type,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire[2:0] T9;
  wire[1:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire T17;
  wire[3:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire[25:0] T22;
  wire[25:0] T23;
  wire[25:0] T24;
  wire T25;
  wire[25:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire[1:0] T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire[1:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire[1:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : 3'h4;
  assign io_out_bits_payload_p_type = T5;
  assign T5 = T13 ? io_in_4_bits_payload_p_type : T6;
  assign T6 = T12 ? T10 : T7;
  assign T7 = T8 ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign T8 = T9[1'h0:1'h0];
  assign T9 = T0;
  assign T10 = T11 ? io_in_3_bits_payload_p_type : io_in_2_bits_payload_p_type;
  assign T11 = T9[1'h0:1'h0];
  assign T12 = T9[1'h1:1'h1];
  assign T13 = T9[2'h2:2'h2];
  assign io_out_bits_payload_master_xact_id = T14;
  assign T14 = T21 ? io_in_4_bits_payload_master_xact_id : T15;
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T17 = T9[1'h0:1'h0];
  assign T18 = T19 ? io_in_3_bits_payload_master_xact_id : io_in_2_bits_payload_master_xact_id;
  assign T19 = T9[1'h0:1'h0];
  assign T20 = T9[1'h1:1'h1];
  assign T21 = T9[2'h2:2'h2];
  assign io_out_bits_payload_addr = T22;
  assign T22 = T29 ? io_in_4_bits_payload_addr : T23;
  assign T23 = T28 ? T26 : T24;
  assign T24 = T25 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T25 = T9[1'h0:1'h0];
  assign T26 = T27 ? io_in_3_bits_payload_addr : io_in_2_bits_payload_addr;
  assign T27 = T9[1'h0:1'h0];
  assign T28 = T9[1'h1:1'h1];
  assign T29 = T9[2'h2:2'h2];
  assign io_out_bits_header_dst = T30;
  assign T30 = T37 ? io_in_4_bits_header_dst : T31;
  assign T31 = T36 ? T34 : T32;
  assign T32 = T33 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T33 = T9[1'h0:1'h0];
  assign T34 = T35 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T35 = T9[1'h0:1'h0];
  assign T36 = T9[1'h1:1'h1];
  assign T37 = T9[2'h2:2'h2];
  assign io_out_bits_header_src = T38;
  assign T38 = T45 ? io_in_4_bits_header_src : T39;
  assign T39 = T44 ? T42 : T40;
  assign T40 = T41 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T41 = T9[1'h0:1'h0];
  assign T42 = T43 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T43 = T9[1'h0:1'h0];
  assign T44 = T9[1'h1:1'h1];
  assign T45 = T9[2'h2:2'h2];
  assign io_out_valid = T46;
  assign T46 = T53 ? io_in_4_valid : T47;
  assign T47 = T52 ? T50 : T48;
  assign T48 = T49 ? io_in_1_valid : io_in_0_valid;
  assign T49 = T9[1'h0:1'h0];
  assign T50 = T51 ? io_in_3_valid : io_in_2_valid;
  assign T51 = T9[1'h0:1'h0];
  assign T52 = T9[1'h1:1'h1];
  assign T53 = T9[2'h2:2'h2];
  assign io_in_0_ready = T54;
  assign T54 = T55 & io_out_ready;
  assign T55 = 1'h1;
  assign io_in_1_ready = T56;
  assign T56 = T57 & io_out_ready;
  assign T57 = T58;
  assign T58 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T59;
  assign T59 = T60 & io_out_ready;
  assign T60 = T61;
  assign T61 = T62 ^ 1'h1;
  assign T62 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T63;
  assign T63 = T64 & io_out_ready;
  assign T64 = T65;
  assign T65 = T66 ^ 1'h1;
  assign T66 = T67 | io_in_2_valid;
  assign T67 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T68;
  assign T68 = T69 & io_out_ready;
  assign T69 = T70;
  assign T70 = T71 ^ 1'h1;
  assign T71 = T72 | io_in_3_valid;
  assign T72 = T73 | io_in_2_valid;
  assign T73 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_13(
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [511:0] io_in_4_bits_payload_data,
    input [3:0] io_in_4_bits_payload_client_xact_id,
    input [3:0] io_in_4_bits_payload_master_xact_id,
    input [3:0] io_in_4_bits_payload_g_type,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [511:0] io_in_3_bits_payload_data,
    input [3:0] io_in_3_bits_payload_client_xact_id,
    input [3:0] io_in_3_bits_payload_master_xact_id,
    input [3:0] io_in_3_bits_payload_g_type,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [511:0] io_in_2_bits_payload_data,
    input [3:0] io_in_2_bits_payload_client_xact_id,
    input [3:0] io_in_2_bits_payload_master_xact_id,
    input [3:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [511:0] io_in_1_bits_payload_data,
    input [3:0] io_in_1_bits_payload_client_xact_id,
    input [3:0] io_in_1_bits_payload_master_xact_id,
    input [3:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [511:0] io_in_0_bits_payload_data,
    input [3:0] io_in_0_bits_payload_client_xact_id,
    input [3:0] io_in_0_bits_payload_master_xact_id,
    input [3:0] io_in_0_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[3:0] io_out_bits_payload_client_xact_id,
    output[3:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire T8;
  wire[2:0] T9;
  wire[3:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire T17;
  wire[3:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire[3:0] T22;
  wire[3:0] T23;
  wire[3:0] T24;
  wire T25;
  wire[3:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire[511:0] T30;
  wire[511:0] T31;
  wire[511:0] T32;
  wire T33;
  wire[511:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire[1:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire[1:0] T46;
  wire[1:0] T47;
  wire[1:0] T48;
  wire T49;
  wire[1:0] T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : 3'h4;
  assign io_out_bits_payload_g_type = T5;
  assign T5 = T13 ? io_in_4_bits_payload_g_type : T6;
  assign T6 = T12 ? T10 : T7;
  assign T7 = T8 ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign T8 = T9[1'h0:1'h0];
  assign T9 = T0;
  assign T10 = T11 ? io_in_3_bits_payload_g_type : io_in_2_bits_payload_g_type;
  assign T11 = T9[1'h0:1'h0];
  assign T12 = T9[1'h1:1'h1];
  assign T13 = T9[2'h2:2'h2];
  assign io_out_bits_payload_master_xact_id = T14;
  assign T14 = T21 ? io_in_4_bits_payload_master_xact_id : T15;
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T17 = T9[1'h0:1'h0];
  assign T18 = T19 ? io_in_3_bits_payload_master_xact_id : io_in_2_bits_payload_master_xact_id;
  assign T19 = T9[1'h0:1'h0];
  assign T20 = T9[1'h1:1'h1];
  assign T21 = T9[2'h2:2'h2];
  assign io_out_bits_payload_client_xact_id = T22;
  assign T22 = T29 ? io_in_4_bits_payload_client_xact_id : T23;
  assign T23 = T28 ? T26 : T24;
  assign T24 = T25 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T25 = T9[1'h0:1'h0];
  assign T26 = T27 ? io_in_3_bits_payload_client_xact_id : io_in_2_bits_payload_client_xact_id;
  assign T27 = T9[1'h0:1'h0];
  assign T28 = T9[1'h1:1'h1];
  assign T29 = T9[2'h2:2'h2];
  assign io_out_bits_payload_data = T30;
  assign T30 = T37 ? io_in_4_bits_payload_data : T31;
  assign T31 = T36 ? T34 : T32;
  assign T32 = T33 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T33 = T9[1'h0:1'h0];
  assign T34 = T35 ? io_in_3_bits_payload_data : io_in_2_bits_payload_data;
  assign T35 = T9[1'h0:1'h0];
  assign T36 = T9[1'h1:1'h1];
  assign T37 = T9[2'h2:2'h2];
  assign io_out_bits_header_dst = T38;
  assign T38 = T45 ? io_in_4_bits_header_dst : T39;
  assign T39 = T44 ? T42 : T40;
  assign T40 = T41 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T41 = T9[1'h0:1'h0];
  assign T42 = T43 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T43 = T9[1'h0:1'h0];
  assign T44 = T9[1'h1:1'h1];
  assign T45 = T9[2'h2:2'h2];
  assign io_out_bits_header_src = T46;
  assign T46 = T53 ? io_in_4_bits_header_src : T47;
  assign T47 = T52 ? T50 : T48;
  assign T48 = T49 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T49 = T9[1'h0:1'h0];
  assign T50 = T51 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T51 = T9[1'h0:1'h0];
  assign T52 = T9[1'h1:1'h1];
  assign T53 = T9[2'h2:2'h2];
  assign io_out_valid = T54;
  assign T54 = T61 ? io_in_4_valid : T55;
  assign T55 = T60 ? T58 : T56;
  assign T56 = T57 ? io_in_1_valid : io_in_0_valid;
  assign T57 = T9[1'h0:1'h0];
  assign T58 = T59 ? io_in_3_valid : io_in_2_valid;
  assign T59 = T9[1'h0:1'h0];
  assign T60 = T9[1'h1:1'h1];
  assign T61 = T9[2'h2:2'h2];
  assign io_in_0_ready = T62;
  assign T62 = T63 & io_out_ready;
  assign T63 = 1'h1;
  assign io_in_1_ready = T64;
  assign T64 = T65 & io_out_ready;
  assign T65 = T66;
  assign T66 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T67;
  assign T67 = T68 & io_out_ready;
  assign T68 = T69;
  assign T69 = T70 ^ 1'h1;
  assign T70 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T71;
  assign T71 = T72 & io_out_ready;
  assign T72 = T73;
  assign T73 = T74 ^ 1'h1;
  assign T74 = T75 | io_in_2_valid;
  assign T75 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T76;
  assign T76 = T77 & io_out_ready;
  assign T77 = T78;
  assign T78 = T79 ^ 1'h1;
  assign T79 = T80 | io_in_3_valid;
  assign T80 = T81 | io_in_2_valid;
  assign T81 = io_in_0_valid | io_in_1_valid;
endmodule

module RRArbiter_3(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr,
    input [3:0] io_in_4_bits_payload_client_xact_id,
    input [511:0] io_in_4_bits_payload_data,
    input [2:0] io_in_4_bits_payload_a_type,
    input [5:0] io_in_4_bits_payload_write_mask,
    input [2:0] io_in_4_bits_payload_subword_addr,
    input [3:0] io_in_4_bits_payload_atomic_opcode,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr,
    input [3:0] io_in_3_bits_payload_client_xact_id,
    input [511:0] io_in_3_bits_payload_data,
    input [2:0] io_in_3_bits_payload_a_type,
    input [5:0] io_in_3_bits_payload_write_mask,
    input [2:0] io_in_3_bits_payload_subword_addr,
    input [3:0] io_in_3_bits_payload_atomic_opcode,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [3:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_a_type,
    input [5:0] io_in_2_bits_payload_write_mask,
    input [2:0] io_in_2_bits_payload_subword_addr,
    input [3:0] io_in_2_bits_payload_atomic_opcode,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [3:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [3:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[3:0] io_out_bits_payload_client_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_a_type,
    output[5:0] io_out_bits_payload_write_mask,
    output[2:0] io_out_bits_payload_subword_addr,
    output[3:0] io_out_bits_payload_atomic_opcode,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;
  reg [2:0] R11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire[3:0] T23;
  wire T24;
  wire[2:0] T25;
  wire[3:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire T33;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire[5:0] T38;
  wire[5:0] T39;
  wire[5:0] T40;
  wire T41;
  wire[5:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire[2:0] T46;
  wire[2:0] T47;
  wire[2:0] T48;
  wire T49;
  wire[2:0] T50;
  wire T51;
  wire T52;
  wire T53;
  wire[511:0] T54;
  wire[511:0] T55;
  wire[511:0] T56;
  wire T57;
  wire[511:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire T65;
  wire[3:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[25:0] T70;
  wire[25:0] T71;
  wire[25:0] T72;
  wire T73;
  wire[25:0] T74;
  wire T75;
  wire T76;
  wire T77;
  wire[1:0] T78;
  wire[1:0] T79;
  wire[1:0] T80;
  wire T81;
  wire[1:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire[1:0] T86;
  wire[1:0] T87;
  wire[1:0] T88;
  wire T89;
  wire[1:0] T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R11 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T19 ? 3'h1 : T2;
  assign T2 = T17 ? 3'h2 : T3;
  assign T3 = T15 ? 3'h3 : T4;
  assign T4 = T9 ? 3'h4 : T5;
  assign T5 = io_in_0_valid ? 3'h0 : T6;
  assign T6 = io_in_1_valid ? 3'h1 : T7;
  assign T7 = io_in_2_valid ? 3'h2 : T8;
  assign T8 = io_in_3_valid ? 3'h3 : 3'h4;
  assign T9 = io_in_4_valid & T10;
  assign T10 = R11 < 3'h4;
  assign T12 = reset ? 3'h0 : T13;
  assign T13 = T14 ? T0 : R11;
  assign T14 = io_out_ready & io_out_valid;
  assign T15 = io_in_3_valid & T16;
  assign T16 = R11 < 3'h3;
  assign T17 = io_in_2_valid & T18;
  assign T18 = R11 < 3'h2;
  assign T19 = io_in_1_valid & T20;
  assign T20 = R11 < 3'h1;
  assign io_out_bits_payload_atomic_opcode = T21;
  assign T21 = T29 ? io_in_4_bits_payload_atomic_opcode : T22;
  assign T22 = T28 ? T26 : T23;
  assign T23 = T24 ? io_in_1_bits_payload_atomic_opcode : io_in_0_bits_payload_atomic_opcode;
  assign T24 = T25[1'h0:1'h0];
  assign T25 = T0;
  assign T26 = T27 ? io_in_3_bits_payload_atomic_opcode : io_in_2_bits_payload_atomic_opcode;
  assign T27 = T25[1'h0:1'h0];
  assign T28 = T25[1'h1:1'h1];
  assign T29 = T25[2'h2:2'h2];
  assign io_out_bits_payload_subword_addr = T30;
  assign T30 = T37 ? io_in_4_bits_payload_subword_addr : T31;
  assign T31 = T36 ? T34 : T32;
  assign T32 = T33 ? io_in_1_bits_payload_subword_addr : io_in_0_bits_payload_subword_addr;
  assign T33 = T25[1'h0:1'h0];
  assign T34 = T35 ? io_in_3_bits_payload_subword_addr : io_in_2_bits_payload_subword_addr;
  assign T35 = T25[1'h0:1'h0];
  assign T36 = T25[1'h1:1'h1];
  assign T37 = T25[2'h2:2'h2];
  assign io_out_bits_payload_write_mask = T38;
  assign T38 = T45 ? io_in_4_bits_payload_write_mask : T39;
  assign T39 = T44 ? T42 : T40;
  assign T40 = T41 ? io_in_1_bits_payload_write_mask : io_in_0_bits_payload_write_mask;
  assign T41 = T25[1'h0:1'h0];
  assign T42 = T43 ? io_in_3_bits_payload_write_mask : io_in_2_bits_payload_write_mask;
  assign T43 = T25[1'h0:1'h0];
  assign T44 = T25[1'h1:1'h1];
  assign T45 = T25[2'h2:2'h2];
  assign io_out_bits_payload_a_type = T46;
  assign T46 = T53 ? io_in_4_bits_payload_a_type : T47;
  assign T47 = T52 ? T50 : T48;
  assign T48 = T49 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T49 = T25[1'h0:1'h0];
  assign T50 = T51 ? io_in_3_bits_payload_a_type : io_in_2_bits_payload_a_type;
  assign T51 = T25[1'h0:1'h0];
  assign T52 = T25[1'h1:1'h1];
  assign T53 = T25[2'h2:2'h2];
  assign io_out_bits_payload_data = T54;
  assign T54 = T61 ? io_in_4_bits_payload_data : T55;
  assign T55 = T60 ? T58 : T56;
  assign T56 = T57 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T57 = T25[1'h0:1'h0];
  assign T58 = T59 ? io_in_3_bits_payload_data : io_in_2_bits_payload_data;
  assign T59 = T25[1'h0:1'h0];
  assign T60 = T25[1'h1:1'h1];
  assign T61 = T25[2'h2:2'h2];
  assign io_out_bits_payload_client_xact_id = T62;
  assign T62 = T69 ? io_in_4_bits_payload_client_xact_id : T63;
  assign T63 = T68 ? T66 : T64;
  assign T64 = T65 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T65 = T25[1'h0:1'h0];
  assign T66 = T67 ? io_in_3_bits_payload_client_xact_id : io_in_2_bits_payload_client_xact_id;
  assign T67 = T25[1'h0:1'h0];
  assign T68 = T25[1'h1:1'h1];
  assign T69 = T25[2'h2:2'h2];
  assign io_out_bits_payload_addr = T70;
  assign T70 = T77 ? io_in_4_bits_payload_addr : T71;
  assign T71 = T76 ? T74 : T72;
  assign T72 = T73 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T73 = T25[1'h0:1'h0];
  assign T74 = T75 ? io_in_3_bits_payload_addr : io_in_2_bits_payload_addr;
  assign T75 = T25[1'h0:1'h0];
  assign T76 = T25[1'h1:1'h1];
  assign T77 = T25[2'h2:2'h2];
  assign io_out_bits_header_dst = T78;
  assign T78 = T85 ? io_in_4_bits_header_dst : T79;
  assign T79 = T84 ? T82 : T80;
  assign T80 = T81 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T81 = T25[1'h0:1'h0];
  assign T82 = T83 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T83 = T25[1'h0:1'h0];
  assign T84 = T25[1'h1:1'h1];
  assign T85 = T25[2'h2:2'h2];
  assign io_out_bits_header_src = T86;
  assign T86 = T93 ? io_in_4_bits_header_src : T87;
  assign T87 = T92 ? T90 : T88;
  assign T88 = T89 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T89 = T25[1'h0:1'h0];
  assign T90 = T91 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T91 = T25[1'h0:1'h0];
  assign T92 = T25[1'h1:1'h1];
  assign T93 = T25[2'h2:2'h2];
  assign io_out_valid = T94;
  assign T94 = T101 ? io_in_4_valid : T95;
  assign T95 = T100 ? T98 : T96;
  assign T96 = T97 ? io_in_1_valid : io_in_0_valid;
  assign T97 = T25[1'h0:1'h0];
  assign T98 = T99 ? io_in_3_valid : io_in_2_valid;
  assign T99 = T25[1'h0:1'h0];
  assign T100 = T25[1'h1:1'h1];
  assign T101 = T25[2'h2:2'h2];
  assign io_in_0_ready = T102;
  assign T102 = T103 & io_out_ready;
  assign T103 = T104;
  assign T104 = T120 | T105;
  assign T105 = T106 ^ 1'h1;
  assign T106 = T109 | T107;
  assign T107 = io_in_4_valid & T108;
  assign T108 = R11 < 3'h4;
  assign T109 = T112 | T110;
  assign T110 = io_in_3_valid & T111;
  assign T111 = R11 < 3'h3;
  assign T112 = T115 | T113;
  assign T113 = io_in_2_valid & T114;
  assign T114 = R11 < 3'h2;
  assign T115 = T118 | T116;
  assign T116 = io_in_1_valid & T117;
  assign T117 = R11 < 3'h1;
  assign T118 = io_in_0_valid & T119;
  assign T119 = R11 < 3'h0;
  assign T120 = R11 < 3'h0;
  assign io_in_1_ready = T121;
  assign T121 = T122 & io_out_ready;
  assign T122 = T123;
  assign T123 = T130 | T124;
  assign T124 = T125 ^ 1'h1;
  assign T125 = T126 | io_in_0_valid;
  assign T126 = T127 | T107;
  assign T127 = T128 | T110;
  assign T128 = T129 | T113;
  assign T129 = T118 | T116;
  assign T130 = T132 & T131;
  assign T131 = R11 < 3'h1;
  assign T132 = T118 ^ 1'h1;
  assign io_in_2_ready = T133;
  assign T133 = T134 & io_out_ready;
  assign T134 = T135;
  assign T135 = T143 | T136;
  assign T136 = T137 ^ 1'h1;
  assign T137 = T138 | io_in_1_valid;
  assign T138 = T139 | io_in_0_valid;
  assign T139 = T140 | T107;
  assign T140 = T141 | T110;
  assign T141 = T142 | T113;
  assign T142 = T118 | T116;
  assign T143 = T145 & T144;
  assign T144 = R11 < 3'h2;
  assign T145 = T146 ^ 1'h1;
  assign T146 = T118 | T116;
  assign io_in_3_ready = T147;
  assign T147 = T148 & io_out_ready;
  assign T148 = T149;
  assign T149 = T158 | T150;
  assign T150 = T151 ^ 1'h1;
  assign T151 = T152 | io_in_2_valid;
  assign T152 = T153 | io_in_1_valid;
  assign T153 = T154 | io_in_0_valid;
  assign T154 = T155 | T107;
  assign T155 = T156 | T110;
  assign T156 = T157 | T113;
  assign T157 = T118 | T116;
  assign T158 = T160 & T159;
  assign T159 = R11 < 3'h3;
  assign T160 = T161 ^ 1'h1;
  assign T161 = T162 | T113;
  assign T162 = T118 | T116;
  assign io_in_4_ready = T163;
  assign T163 = T164 & io_out_ready;
  assign T164 = T165;
  assign T165 = T175 | T166;
  assign T166 = T167 ^ 1'h1;
  assign T167 = T168 | io_in_3_valid;
  assign T168 = T169 | io_in_2_valid;
  assign T169 = T170 | io_in_1_valid;
  assign T170 = T171 | io_in_0_valid;
  assign T171 = T172 | T107;
  assign T172 = T173 | T110;
  assign T173 = T174 | T113;
  assign T174 = T118 | T116;
  assign T175 = T177 & T176;
  assign T176 = R11 < 3'h4;
  assign T177 = T178 ^ 1'h1;
  assign T178 = T179 | T110;
  assign T179 = T180 | T113;
  assign T180 = T118 | T116;

  always @(posedge clk) begin
    if(reset) begin
      R11 <= 3'h0;
    end else if(T14) begin
      R11 <= T0;
    end
  end
endmodule

module RRArbiter_4(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [3:0] io_in_4_bits_payload_master_xact_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [3:0] io_in_3_bits_payload_master_xact_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [3:0] io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [3:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [3:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[3:0] io_out_bits_payload_master_xact_id,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire T9;
  wire T10;
  reg [2:0] R11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire[3:0] T23;
  wire T24;
  wire[2:0] T25;
  wire[3:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire[1:0] T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire[1:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire[1:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R11 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T19 ? 3'h1 : T2;
  assign T2 = T17 ? 3'h2 : T3;
  assign T3 = T15 ? 3'h3 : T4;
  assign T4 = T9 ? 3'h4 : T5;
  assign T5 = io_in_0_valid ? 3'h0 : T6;
  assign T6 = io_in_1_valid ? 3'h1 : T7;
  assign T7 = io_in_2_valid ? 3'h2 : T8;
  assign T8 = io_in_3_valid ? 3'h3 : 3'h4;
  assign T9 = io_in_4_valid & T10;
  assign T10 = R11 < 3'h4;
  assign T12 = reset ? 3'h0 : T13;
  assign T13 = T14 ? T0 : R11;
  assign T14 = io_out_ready & io_out_valid;
  assign T15 = io_in_3_valid & T16;
  assign T16 = R11 < 3'h3;
  assign T17 = io_in_2_valid & T18;
  assign T18 = R11 < 3'h2;
  assign T19 = io_in_1_valid & T20;
  assign T20 = R11 < 3'h1;
  assign io_out_bits_payload_master_xact_id = T21;
  assign T21 = T29 ? io_in_4_bits_payload_master_xact_id : T22;
  assign T22 = T28 ? T26 : T23;
  assign T23 = T24 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T24 = T25[1'h0:1'h0];
  assign T25 = T0;
  assign T26 = T27 ? io_in_3_bits_payload_master_xact_id : io_in_2_bits_payload_master_xact_id;
  assign T27 = T25[1'h0:1'h0];
  assign T28 = T25[1'h1:1'h1];
  assign T29 = T25[2'h2:2'h2];
  assign io_out_bits_header_dst = T30;
  assign T30 = T37 ? io_in_4_bits_header_dst : T31;
  assign T31 = T36 ? T34 : T32;
  assign T32 = T33 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T33 = T25[1'h0:1'h0];
  assign T34 = T35 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T35 = T25[1'h0:1'h0];
  assign T36 = T25[1'h1:1'h1];
  assign T37 = T25[2'h2:2'h2];
  assign io_out_bits_header_src = T38;
  assign T38 = T45 ? io_in_4_bits_header_src : T39;
  assign T39 = T44 ? T42 : T40;
  assign T40 = T41 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T41 = T25[1'h0:1'h0];
  assign T42 = T43 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T43 = T25[1'h0:1'h0];
  assign T44 = T25[1'h1:1'h1];
  assign T45 = T25[2'h2:2'h2];
  assign io_out_valid = T46;
  assign T46 = T53 ? io_in_4_valid : T47;
  assign T47 = T52 ? T50 : T48;
  assign T48 = T49 ? io_in_1_valid : io_in_0_valid;
  assign T49 = T25[1'h0:1'h0];
  assign T50 = T51 ? io_in_3_valid : io_in_2_valid;
  assign T51 = T25[1'h0:1'h0];
  assign T52 = T25[1'h1:1'h1];
  assign T53 = T25[2'h2:2'h2];
  assign io_in_0_ready = T54;
  assign T54 = T55 & io_out_ready;
  assign T55 = T56;
  assign T56 = T72 | T57;
  assign T57 = T58 ^ 1'h1;
  assign T58 = T61 | T59;
  assign T59 = io_in_4_valid & T60;
  assign T60 = R11 < 3'h4;
  assign T61 = T64 | T62;
  assign T62 = io_in_3_valid & T63;
  assign T63 = R11 < 3'h3;
  assign T64 = T67 | T65;
  assign T65 = io_in_2_valid & T66;
  assign T66 = R11 < 3'h2;
  assign T67 = T70 | T68;
  assign T68 = io_in_1_valid & T69;
  assign T69 = R11 < 3'h1;
  assign T70 = io_in_0_valid & T71;
  assign T71 = R11 < 3'h0;
  assign T72 = R11 < 3'h0;
  assign io_in_1_ready = T73;
  assign T73 = T74 & io_out_ready;
  assign T74 = T75;
  assign T75 = T82 | T76;
  assign T76 = T77 ^ 1'h1;
  assign T77 = T78 | io_in_0_valid;
  assign T78 = T79 | T59;
  assign T79 = T80 | T62;
  assign T80 = T81 | T65;
  assign T81 = T70 | T68;
  assign T82 = T84 & T83;
  assign T83 = R11 < 3'h1;
  assign T84 = T70 ^ 1'h1;
  assign io_in_2_ready = T85;
  assign T85 = T86 & io_out_ready;
  assign T86 = T87;
  assign T87 = T95 | T88;
  assign T88 = T89 ^ 1'h1;
  assign T89 = T90 | io_in_1_valid;
  assign T90 = T91 | io_in_0_valid;
  assign T91 = T92 | T59;
  assign T92 = T93 | T62;
  assign T93 = T94 | T65;
  assign T94 = T70 | T68;
  assign T95 = T97 & T96;
  assign T96 = R11 < 3'h2;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T70 | T68;
  assign io_in_3_ready = T99;
  assign T99 = T100 & io_out_ready;
  assign T100 = T101;
  assign T101 = T110 | T102;
  assign T102 = T103 ^ 1'h1;
  assign T103 = T104 | io_in_2_valid;
  assign T104 = T105 | io_in_1_valid;
  assign T105 = T106 | io_in_0_valid;
  assign T106 = T107 | T59;
  assign T107 = T108 | T62;
  assign T108 = T109 | T65;
  assign T109 = T70 | T68;
  assign T110 = T112 & T111;
  assign T111 = R11 < 3'h3;
  assign T112 = T113 ^ 1'h1;
  assign T113 = T114 | T65;
  assign T114 = T70 | T68;
  assign io_in_4_ready = T115;
  assign T115 = T116 & io_out_ready;
  assign T116 = T117;
  assign T117 = T127 | T118;
  assign T118 = T119 ^ 1'h1;
  assign T119 = T120 | io_in_3_valid;
  assign T120 = T121 | io_in_2_valid;
  assign T121 = T122 | io_in_1_valid;
  assign T122 = T123 | io_in_0_valid;
  assign T123 = T124 | T59;
  assign T124 = T125 | T62;
  assign T125 = T126 | T65;
  assign T126 = T70 | T68;
  assign T127 = T129 & T128;
  assign T128 = R11 < 3'h4;
  assign T129 = T130 ^ 1'h1;
  assign T130 = T131 | T62;
  assign T131 = T132 | T65;
  assign T132 = T70 | T68;

  always @(posedge clk) begin
    if(reset) begin
      R11 <= 3'h0;
    end else if(T14) begin
      R11 <= T0;
    end
  end
endmodule

module UncachedTileLinkIOArbiterThatPassesId(input clk, input reset,
    output io_in_4_acquire_ready,
    input  io_in_4_acquire_valid,
    input [1:0] io_in_4_acquire_bits_header_src,
    input [1:0] io_in_4_acquire_bits_header_dst,
    input [25:0] io_in_4_acquire_bits_payload_addr,
    input [3:0] io_in_4_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_4_acquire_bits_payload_data,
    input [2:0] io_in_4_acquire_bits_payload_a_type,
    input [5:0] io_in_4_acquire_bits_payload_write_mask,
    input [2:0] io_in_4_acquire_bits_payload_subword_addr,
    input [3:0] io_in_4_acquire_bits_payload_atomic_opcode,
    input  io_in_4_grant_ready,
    output io_in_4_grant_valid,
    output[1:0] io_in_4_grant_bits_header_src,
    output[1:0] io_in_4_grant_bits_header_dst,
    output[511:0] io_in_4_grant_bits_payload_data,
    output[3:0] io_in_4_grant_bits_payload_client_xact_id,
    output[3:0] io_in_4_grant_bits_payload_master_xact_id,
    output[3:0] io_in_4_grant_bits_payload_g_type,
    output io_in_4_finish_ready,
    input  io_in_4_finish_valid,
    input [1:0] io_in_4_finish_bits_header_src,
    input [1:0] io_in_4_finish_bits_header_dst,
    input [3:0] io_in_4_finish_bits_payload_master_xact_id,
    output io_in_3_acquire_ready,
    input  io_in_3_acquire_valid,
    input [1:0] io_in_3_acquire_bits_header_src,
    input [1:0] io_in_3_acquire_bits_header_dst,
    input [25:0] io_in_3_acquire_bits_payload_addr,
    input [3:0] io_in_3_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_3_acquire_bits_payload_data,
    input [2:0] io_in_3_acquire_bits_payload_a_type,
    input [5:0] io_in_3_acquire_bits_payload_write_mask,
    input [2:0] io_in_3_acquire_bits_payload_subword_addr,
    input [3:0] io_in_3_acquire_bits_payload_atomic_opcode,
    input  io_in_3_grant_ready,
    output io_in_3_grant_valid,
    output[1:0] io_in_3_grant_bits_header_src,
    output[1:0] io_in_3_grant_bits_header_dst,
    output[511:0] io_in_3_grant_bits_payload_data,
    output[3:0] io_in_3_grant_bits_payload_client_xact_id,
    output[3:0] io_in_3_grant_bits_payload_master_xact_id,
    output[3:0] io_in_3_grant_bits_payload_g_type,
    output io_in_3_finish_ready,
    input  io_in_3_finish_valid,
    input [1:0] io_in_3_finish_bits_header_src,
    input [1:0] io_in_3_finish_bits_header_dst,
    input [3:0] io_in_3_finish_bits_payload_master_xact_id,
    output io_in_2_acquire_ready,
    input  io_in_2_acquire_valid,
    input [1:0] io_in_2_acquire_bits_header_src,
    input [1:0] io_in_2_acquire_bits_header_dst,
    input [25:0] io_in_2_acquire_bits_payload_addr,
    input [3:0] io_in_2_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_2_acquire_bits_payload_data,
    input [2:0] io_in_2_acquire_bits_payload_a_type,
    input [5:0] io_in_2_acquire_bits_payload_write_mask,
    input [2:0] io_in_2_acquire_bits_payload_subword_addr,
    input [3:0] io_in_2_acquire_bits_payload_atomic_opcode,
    input  io_in_2_grant_ready,
    output io_in_2_grant_valid,
    output[1:0] io_in_2_grant_bits_header_src,
    output[1:0] io_in_2_grant_bits_header_dst,
    output[511:0] io_in_2_grant_bits_payload_data,
    output[3:0] io_in_2_grant_bits_payload_client_xact_id,
    output[3:0] io_in_2_grant_bits_payload_master_xact_id,
    output[3:0] io_in_2_grant_bits_payload_g_type,
    output io_in_2_finish_ready,
    input  io_in_2_finish_valid,
    input [1:0] io_in_2_finish_bits_header_src,
    input [1:0] io_in_2_finish_bits_header_dst,
    input [3:0] io_in_2_finish_bits_payload_master_xact_id,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [1:0] io_in_1_acquire_bits_header_src,
    input [1:0] io_in_1_acquire_bits_header_dst,
    input [25:0] io_in_1_acquire_bits_payload_addr,
    input [3:0] io_in_1_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_1_acquire_bits_payload_data,
    input [2:0] io_in_1_acquire_bits_payload_a_type,
    input [5:0] io_in_1_acquire_bits_payload_write_mask,
    input [2:0] io_in_1_acquire_bits_payload_subword_addr,
    input [3:0] io_in_1_acquire_bits_payload_atomic_opcode,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_header_src,
    output[1:0] io_in_1_grant_bits_header_dst,
    output[511:0] io_in_1_grant_bits_payload_data,
    output[3:0] io_in_1_grant_bits_payload_client_xact_id,
    output[3:0] io_in_1_grant_bits_payload_master_xact_id,
    output[3:0] io_in_1_grant_bits_payload_g_type,
    output io_in_1_finish_ready,
    input  io_in_1_finish_valid,
    input [1:0] io_in_1_finish_bits_header_src,
    input [1:0] io_in_1_finish_bits_header_dst,
    input [3:0] io_in_1_finish_bits_payload_master_xact_id,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [1:0] io_in_0_acquire_bits_header_src,
    input [1:0] io_in_0_acquire_bits_header_dst,
    input [25:0] io_in_0_acquire_bits_payload_addr,
    input [3:0] io_in_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_0_acquire_bits_payload_data,
    input [2:0] io_in_0_acquire_bits_payload_a_type,
    input [5:0] io_in_0_acquire_bits_payload_write_mask,
    input [2:0] io_in_0_acquire_bits_payload_subword_addr,
    input [3:0] io_in_0_acquire_bits_payload_atomic_opcode,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_header_src,
    output[1:0] io_in_0_grant_bits_header_dst,
    output[511:0] io_in_0_grant_bits_payload_data,
    output[3:0] io_in_0_grant_bits_payload_client_xact_id,
    output[3:0] io_in_0_grant_bits_payload_master_xact_id,
    output[3:0] io_in_0_grant_bits_payload_g_type,
    output io_in_0_finish_ready,
    input  io_in_0_finish_valid,
    input [1:0] io_in_0_finish_bits_header_src,
    input [1:0] io_in_0_finish_bits_header_dst,
    input [3:0] io_in_0_finish_bits_payload_master_xact_id,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[1:0] io_out_acquire_bits_header_src,
    output[1:0] io_out_acquire_bits_header_dst,
    output[25:0] io_out_acquire_bits_payload_addr,
    output[3:0] io_out_acquire_bits_payload_client_xact_id,
    output[511:0] io_out_acquire_bits_payload_data,
    output[2:0] io_out_acquire_bits_payload_a_type,
    output[5:0] io_out_acquire_bits_payload_write_mask,
    output[2:0] io_out_acquire_bits_payload_subword_addr,
    output[3:0] io_out_acquire_bits_payload_atomic_opcode,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_header_src,
    input [1:0] io_out_grant_bits_header_dst,
    input [511:0] io_out_grant_bits_payload_data,
    input [3:0] io_out_grant_bits_payload_client_xact_id,
    input [3:0] io_out_grant_bits_payload_master_xact_id,
    input [3:0] io_out_grant_bits_payload_g_type,
    input  io_out_finish_ready,
    output io_out_finish_valid,
    output[1:0] io_out_finish_bits_header_src,
    output[1:0] io_out_finish_bits_header_dst,
    output[3:0] io_out_finish_bits_payload_master_xact_id
);

  wire[3:0] RRArbiter_1_io_out_bits_payload_master_xact_id;
  wire[1:0] RRArbiter_1_io_out_bits_header_dst;
  wire[1:0] RRArbiter_1_io_out_bits_header_src;
  wire RRArbiter_1_io_out_valid;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire[3:0] RRArbiter_0_io_out_bits_payload_atomic_opcode;
  wire[2:0] RRArbiter_0_io_out_bits_payload_subword_addr;
  wire[5:0] RRArbiter_0_io_out_bits_payload_write_mask;
  wire[2:0] RRArbiter_0_io_out_bits_payload_a_type;
  wire[511:0] RRArbiter_0_io_out_bits_payload_data;
  wire[3:0] RRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[25:0] RRArbiter_0_io_out_bits_payload_addr;
  wire[1:0] RRArbiter_0_io_out_bits_header_dst;
  wire[1:0] RRArbiter_0_io_out_bits_header_src;
  wire RRArbiter_0_io_out_valid;
  wire RRArbiter_1_io_in_0_ready;
  wire T10;
  wire RRArbiter_0_io_in_0_ready;
  wire RRArbiter_1_io_in_1_ready;
  wire T11;
  wire RRArbiter_0_io_in_1_ready;
  wire RRArbiter_1_io_in_2_ready;
  wire T12;
  wire RRArbiter_0_io_in_2_ready;
  wire RRArbiter_1_io_in_3_ready;
  wire T13;
  wire RRArbiter_0_io_in_3_ready;
  wire RRArbiter_1_io_in_4_ready;
  wire T14;
  wire RRArbiter_0_io_in_4_ready;


  assign io_out_finish_bits_payload_master_xact_id = RRArbiter_1_io_out_bits_payload_master_xact_id;
  assign io_out_finish_bits_header_dst = RRArbiter_1_io_out_bits_header_dst;
  assign io_out_finish_bits_header_src = RRArbiter_1_io_out_bits_header_src;
  assign io_out_finish_valid = RRArbiter_1_io_out_valid;
  assign io_out_grant_ready = T0;
  assign T0 = T9 ? io_in_4_grant_ready : T1;
  assign T1 = T8 ? io_in_3_grant_ready : T2;
  assign T2 = T7 ? io_in_2_grant_ready : T3;
  assign T3 = T6 ? io_in_1_grant_ready : T4;
  assign T4 = T5 ? io_in_0_grant_ready : 1'h0;
  assign T5 = io_out_grant_bits_payload_client_xact_id == 4'h0;
  assign T6 = io_out_grant_bits_payload_client_xact_id == 4'h1;
  assign T7 = io_out_grant_bits_payload_client_xact_id == 4'h2;
  assign T8 = io_out_grant_bits_payload_client_xact_id == 4'h3;
  assign T9 = io_out_grant_bits_payload_client_xact_id == 4'h4;
  assign io_out_acquire_bits_payload_atomic_opcode = RRArbiter_0_io_out_bits_payload_atomic_opcode;
  assign io_out_acquire_bits_payload_subword_addr = RRArbiter_0_io_out_bits_payload_subword_addr;
  assign io_out_acquire_bits_payload_write_mask = RRArbiter_0_io_out_bits_payload_write_mask;
  assign io_out_acquire_bits_payload_a_type = RRArbiter_0_io_out_bits_payload_a_type;
  assign io_out_acquire_bits_payload_data = RRArbiter_0_io_out_bits_payload_data;
  assign io_out_acquire_bits_payload_client_xact_id = RRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_acquire_bits_payload_addr = RRArbiter_0_io_out_bits_payload_addr;
  assign io_out_acquire_bits_header_dst = RRArbiter_0_io_out_bits_header_dst;
  assign io_out_acquire_bits_header_src = RRArbiter_0_io_out_bits_header_src;
  assign io_out_acquire_valid = RRArbiter_0_io_out_valid;
  assign io_in_0_finish_ready = RRArbiter_1_io_in_0_ready;
  assign io_in_0_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_0_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_0_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_0_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_0_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_0_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_0_grant_valid = T10;
  assign T10 = T5 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = RRArbiter_0_io_in_0_ready;
  assign io_in_1_finish_ready = RRArbiter_1_io_in_1_ready;
  assign io_in_1_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_1_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_1_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_1_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_1_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_1_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_1_grant_valid = T11;
  assign T11 = T6 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = RRArbiter_0_io_in_1_ready;
  assign io_in_2_finish_ready = RRArbiter_1_io_in_2_ready;
  assign io_in_2_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_2_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_2_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_2_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_2_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_2_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_2_grant_valid = T12;
  assign T12 = T7 ? io_out_grant_valid : 1'h0;
  assign io_in_2_acquire_ready = RRArbiter_0_io_in_2_ready;
  assign io_in_3_finish_ready = RRArbiter_1_io_in_3_ready;
  assign io_in_3_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_3_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_3_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_3_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_3_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_3_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_3_grant_valid = T13;
  assign T13 = T8 ? io_out_grant_valid : 1'h0;
  assign io_in_3_acquire_ready = RRArbiter_0_io_in_3_ready;
  assign io_in_4_finish_ready = RRArbiter_1_io_in_4_ready;
  assign io_in_4_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_4_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_4_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_4_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_4_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_4_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_4_grant_valid = T14;
  assign T14 = T9 ? io_out_grant_valid : 1'h0;
  assign io_in_4_acquire_ready = RRArbiter_0_io_in_4_ready;
  RRArbiter_3 RRArbiter_0(.clk(clk), .reset(reset),
       .io_in_4_ready( RRArbiter_0_io_in_4_ready ),
       .io_in_4_valid( io_in_4_acquire_valid ),
       .io_in_4_bits_header_src( io_in_4_acquire_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_acquire_bits_header_dst ),
       .io_in_4_bits_payload_addr( io_in_4_acquire_bits_payload_addr ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_acquire_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_data( io_in_4_acquire_bits_payload_data ),
       .io_in_4_bits_payload_a_type( io_in_4_acquire_bits_payload_a_type ),
       .io_in_4_bits_payload_write_mask( io_in_4_acquire_bits_payload_write_mask ),
       .io_in_4_bits_payload_subword_addr( io_in_4_acquire_bits_payload_subword_addr ),
       .io_in_4_bits_payload_atomic_opcode( io_in_4_acquire_bits_payload_atomic_opcode ),
       .io_in_3_ready( RRArbiter_0_io_in_3_ready ),
       .io_in_3_valid( io_in_3_acquire_valid ),
       .io_in_3_bits_header_src( io_in_3_acquire_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_acquire_bits_header_dst ),
       .io_in_3_bits_payload_addr( io_in_3_acquire_bits_payload_addr ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_acquire_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_data( io_in_3_acquire_bits_payload_data ),
       .io_in_3_bits_payload_a_type( io_in_3_acquire_bits_payload_a_type ),
       .io_in_3_bits_payload_write_mask( io_in_3_acquire_bits_payload_write_mask ),
       .io_in_3_bits_payload_subword_addr( io_in_3_acquire_bits_payload_subword_addr ),
       .io_in_3_bits_payload_atomic_opcode( io_in_3_acquire_bits_payload_atomic_opcode ),
       .io_in_2_ready( RRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( io_in_2_acquire_valid ),
       .io_in_2_bits_header_src( io_in_2_acquire_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_acquire_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_acquire_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_acquire_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_acquire_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_acquire_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_acquire_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_acquire_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_acquire_bits_payload_atomic_opcode ),
       .io_in_1_ready( RRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_header_src( io_in_1_acquire_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_acquire_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_acquire_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_acquire_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_acquire_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_acquire_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_acquire_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_acquire_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_acquire_bits_payload_atomic_opcode ),
       .io_in_0_ready( RRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_header_src( io_in_0_acquire_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_acquire_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_acquire_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_acquire_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_acquire_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_acquire_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_acquire_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_acquire_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_acquire_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( RRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( RRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( RRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( RRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( RRArbiter_0_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( RRArbiter_0_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( RRArbiter_0_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( RRArbiter_0_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  RRArbiter_4 RRArbiter_1(.clk(clk), .reset(reset),
       .io_in_4_ready( RRArbiter_1_io_in_4_ready ),
       .io_in_4_valid( io_in_4_finish_valid ),
       .io_in_4_bits_header_src( io_in_4_finish_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_finish_bits_header_dst ),
       .io_in_4_bits_payload_master_xact_id( io_in_4_finish_bits_payload_master_xact_id ),
       .io_in_3_ready( RRArbiter_1_io_in_3_ready ),
       .io_in_3_valid( io_in_3_finish_valid ),
       .io_in_3_bits_header_src( io_in_3_finish_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_finish_bits_header_dst ),
       .io_in_3_bits_payload_master_xact_id( io_in_3_finish_bits_payload_master_xact_id ),
       .io_in_2_ready( RRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( io_in_2_finish_valid ),
       .io_in_2_bits_header_src( io_in_2_finish_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_finish_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_finish_bits_payload_master_xact_id ),
       .io_in_1_ready( RRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( io_in_1_finish_valid ),
       .io_in_1_bits_header_src( io_in_1_finish_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_finish_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_finish_bits_payload_master_xact_id ),
       .io_in_0_ready( RRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( io_in_0_finish_valid ),
       .io_in_0_bits_header_src( io_in_0_finish_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_finish_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_finish_bits_payload_master_xact_id ),
       .io_out_ready( io_out_finish_ready ),
       .io_out_valid( RRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( RRArbiter_1_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
endmodule

module L2CoherenceAgent(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [3:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[3:0] io_inner_grant_bits_payload_client_xact_id,
    output[3:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [3:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[3:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [3:0] io_inner_release_bits_payload_client_xact_id,
    input [3:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    output[1:0] io_outer_acquire_bits_header_dst,
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[3:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [3:0] io_outer_grant_bits_payload_client_xact_id,
    input [3:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    output io_outer_finish_valid,
    output[1:0] io_outer_finish_bits_header_src,
    output[1:0] io_outer_finish_bits_header_dst,
    output[3:0] io_outer_finish_bits_payload_master_xact_id,
    input  io_incoherent_1,
    input  io_incoherent_0
);

  wire VoluntaryReleaseTracker_io_outer_grant_ready;
  wire[3:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_atomic_opcode;
  wire[2:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subword_addr;
  wire[5:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type;
  wire[511:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data;
  wire[3:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id;
  wire[25:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr;
  wire[1:0] VoluntaryReleaseTracker_io_outer_acquire_bits_header_src;
  wire VoluntaryReleaseTracker_io_outer_acquire_valid;
  wire AcquireTracker_0_io_outer_grant_ready;
  wire[3:0] AcquireTracker_0_io_outer_acquire_bits_payload_atomic_opcode;
  wire[2:0] AcquireTracker_0_io_outer_acquire_bits_payload_subword_addr;
  wire[5:0] AcquireTracker_0_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_0_io_outer_acquire_bits_payload_a_type;
  wire[511:0] AcquireTracker_0_io_outer_acquire_bits_payload_data;
  wire[3:0] AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id;
  wire[25:0] AcquireTracker_0_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_0_io_outer_acquire_bits_header_src;
  wire AcquireTracker_0_io_outer_acquire_valid;
  wire AcquireTracker_1_io_outer_grant_ready;
  wire[3:0] AcquireTracker_1_io_outer_acquire_bits_payload_atomic_opcode;
  wire[2:0] AcquireTracker_1_io_outer_acquire_bits_payload_subword_addr;
  wire[5:0] AcquireTracker_1_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_1_io_outer_acquire_bits_payload_a_type;
  wire[511:0] AcquireTracker_1_io_outer_acquire_bits_payload_data;
  wire[3:0] AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id;
  wire[25:0] AcquireTracker_1_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_1_io_outer_acquire_bits_header_src;
  wire AcquireTracker_1_io_outer_acquire_valid;
  wire AcquireTracker_2_io_outer_grant_ready;
  wire[3:0] AcquireTracker_2_io_outer_acquire_bits_payload_atomic_opcode;
  wire[2:0] AcquireTracker_2_io_outer_acquire_bits_payload_subword_addr;
  wire[5:0] AcquireTracker_2_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_2_io_outer_acquire_bits_payload_a_type;
  wire[511:0] AcquireTracker_2_io_outer_acquire_bits_payload_data;
  wire[3:0] AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id;
  wire[25:0] AcquireTracker_2_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_2_io_outer_acquire_bits_header_src;
  wire AcquireTracker_2_io_outer_acquire_valid;
  wire AcquireTracker_3_io_outer_grant_ready;
  wire[3:0] AcquireTracker_3_io_outer_acquire_bits_payload_atomic_opcode;
  wire[2:0] AcquireTracker_3_io_outer_acquire_bits_payload_subword_addr;
  wire[5:0] AcquireTracker_3_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_3_io_outer_acquire_bits_payload_a_type;
  wire[511:0] AcquireTracker_3_io_outer_acquire_bits_payload_data;
  wire[3:0] AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id;
  wire[25:0] AcquireTracker_3_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_3_io_outer_acquire_bits_header_src;
  wire AcquireTracker_3_io_outer_acquire_valid;
  wire[3:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type;
  wire[3:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id;
  wire[511:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_data;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_header_dst;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_header_src;
  wire VoluntaryReleaseTracker_io_inner_grant_valid;
  wire[3:0] AcquireTracker_0_io_inner_grant_bits_payload_g_type;
  wire[3:0] AcquireTracker_0_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_0_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_header_dst;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_header_src;
  wire AcquireTracker_0_io_inner_grant_valid;
  wire[3:0] AcquireTracker_1_io_inner_grant_bits_payload_g_type;
  wire[3:0] AcquireTracker_1_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_1_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_header_dst;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_header_src;
  wire AcquireTracker_1_io_inner_grant_valid;
  wire[3:0] AcquireTracker_2_io_inner_grant_bits_payload_g_type;
  wire[3:0] AcquireTracker_2_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_2_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_header_dst;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_header_src;
  wire AcquireTracker_2_io_inner_grant_valid;
  wire[3:0] AcquireTracker_3_io_inner_grant_bits_payload_g_type;
  wire[3:0] AcquireTracker_3_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_3_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_header_dst;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_header_src;
  wire AcquireTracker_3_io_inner_grant_valid;
  wire VoluntaryReleaseTracker_io_inner_probe_valid;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_payload_p_type;
  wire[3:0] AcquireTracker_0_io_inner_probe_bits_payload_master_xact_id;
  wire[25:0] AcquireTracker_0_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_header_dst;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_header_src;
  wire AcquireTracker_0_io_inner_probe_valid;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_payload_p_type;
  wire[3:0] AcquireTracker_1_io_inner_probe_bits_payload_master_xact_id;
  wire[25:0] AcquireTracker_1_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_header_dst;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_header_src;
  wire AcquireTracker_1_io_inner_probe_valid;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_payload_p_type;
  wire[3:0] AcquireTracker_2_io_inner_probe_bits_payload_master_xact_id;
  wire[25:0] AcquireTracker_2_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_header_dst;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_header_src;
  wire AcquireTracker_2_io_inner_probe_valid;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_payload_p_type;
  wire[3:0] AcquireTracker_3_io_inner_probe_bits_payload_master_xact_id;
  wire[25:0] AcquireTracker_3_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_header_dst;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_header_src;
  wire AcquireTracker_3_io_inner_probe_valid;
  wire T0;
  wire T1;
  wire block_acquires;
  wire AcquireTracker_3_io_has_acquire_conflict;
  wire T2;
  wire AcquireTracker_2_io_has_acquire_conflict;
  wire T3;
  wire AcquireTracker_1_io_has_acquire_conflict;
  wire T4;
  wire AcquireTracker_0_io_has_acquire_conflict;
  wire VoluntaryReleaseTracker_io_has_acquire_conflict;
  wire VoluntaryReleaseTracker_io_inner_acquire_ready;
  wire AcquireTracker_0_io_inner_acquire_ready;
  wire AcquireTracker_1_io_inner_acquire_ready;
  wire AcquireTracker_2_io_inner_acquire_ready;
  wire AcquireTracker_3_io_inner_acquire_ready;
  wire[1:0] T5;
  wire[1:0] T6;
  wire outer_arb_io_in_4_finish_ready;
  wire[3:0] outer_arb_io_in_4_grant_bits_payload_g_type;
  wire[3:0] outer_arb_io_in_4_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_4_grant_bits_payload_client_xact_id;
  wire[511:0] outer_arb_io_in_4_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_4_grant_bits_header_dst;
  wire[1:0] outer_arb_io_in_4_grant_bits_header_src;
  wire outer_arb_io_in_4_grant_valid;
  wire outer_arb_io_in_4_acquire_ready;
  wire T7;
  wire T8;
  wire[3:0] release_idx;
  wire voluntary;
  wire probe_arb_io_in_4_ready;
  wire grant_arb_io_in_4_ready;
  wire alloc_arb_io_in_4_ready;
  wire[1:0] T9;
  wire outer_arb_io_in_3_finish_ready;
  wire[3:0] outer_arb_io_in_3_grant_bits_payload_g_type;
  wire[3:0] outer_arb_io_in_3_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_3_grant_bits_payload_client_xact_id;
  wire[511:0] outer_arb_io_in_3_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_3_grant_bits_header_dst;
  wire[1:0] outer_arb_io_in_3_grant_bits_header_src;
  wire outer_arb_io_in_3_grant_valid;
  wire outer_arb_io_in_3_acquire_ready;
  wire T10;
  wire T11;
  wire probe_arb_io_in_3_ready;
  wire grant_arb_io_in_3_ready;
  wire alloc_arb_io_in_3_ready;
  wire[1:0] T12;
  wire outer_arb_io_in_2_finish_ready;
  wire[3:0] outer_arb_io_in_2_grant_bits_payload_g_type;
  wire[3:0] outer_arb_io_in_2_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_2_grant_bits_payload_client_xact_id;
  wire[511:0] outer_arb_io_in_2_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_2_grant_bits_header_dst;
  wire[1:0] outer_arb_io_in_2_grant_bits_header_src;
  wire outer_arb_io_in_2_grant_valid;
  wire outer_arb_io_in_2_acquire_ready;
  wire T13;
  wire T14;
  wire probe_arb_io_in_2_ready;
  wire grant_arb_io_in_2_ready;
  wire alloc_arb_io_in_2_ready;
  wire[1:0] T15;
  wire outer_arb_io_in_1_finish_ready;
  wire[3:0] outer_arb_io_in_1_grant_bits_payload_g_type;
  wire[3:0] outer_arb_io_in_1_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_1_grant_bits_payload_client_xact_id;
  wire[511:0] outer_arb_io_in_1_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_1_grant_bits_header_dst;
  wire[1:0] outer_arb_io_in_1_grant_bits_header_src;
  wire outer_arb_io_in_1_grant_valid;
  wire outer_arb_io_in_1_acquire_ready;
  wire T16;
  wire T17;
  wire probe_arb_io_in_1_ready;
  wire grant_arb_io_in_1_ready;
  wire alloc_arb_io_in_1_ready;
  wire[1:0] T18;
  wire outer_arb_io_in_0_finish_ready;
  wire[3:0] outer_arb_io_in_0_grant_bits_payload_g_type;
  wire[3:0] outer_arb_io_in_0_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_0_grant_bits_payload_client_xact_id;
  wire[511:0] outer_arb_io_in_0_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_0_grant_bits_header_dst;
  wire[1:0] outer_arb_io_in_0_grant_bits_header_src;
  wire outer_arb_io_in_0_grant_valid;
  wire outer_arb_io_in_0_acquire_ready;
  wire T19;
  wire T20;
  wire probe_arb_io_in_0_ready;
  wire grant_arb_io_in_0_ready;
  wire alloc_arb_io_in_0_ready;
  wire[3:0] outer_arb_io_out_finish_bits_payload_master_xact_id;
  wire[1:0] outer_arb_io_out_finish_bits_header_dst;
  wire[1:0] outer_arb_io_out_finish_bits_header_src;
  wire outer_arb_io_out_finish_valid;
  wire outer_arb_io_out_grant_ready;
  wire[3:0] outer_arb_io_out_acquire_bits_payload_atomic_opcode;
  wire[2:0] outer_arb_io_out_acquire_bits_payload_subword_addr;
  wire[5:0] outer_arb_io_out_acquire_bits_payload_write_mask;
  wire[2:0] outer_arb_io_out_acquire_bits_payload_a_type;
  wire[511:0] outer_arb_io_out_acquire_bits_payload_data;
  wire[3:0] outer_arb_io_out_acquire_bits_payload_client_xact_id;
  wire[25:0] outer_arb_io_out_acquire_bits_payload_addr;
  wire[1:0] outer_arb_io_out_acquire_bits_header_dst;
  wire[1:0] outer_arb_io_out_acquire_bits_header_src;
  wire outer_arb_io_out_acquire_valid;
  wire T21;
  wire T22;
  wire T23;
  wire VoluntaryReleaseTracker_io_inner_release_ready;
  wire AcquireTracker_0_io_inner_release_ready;
  wire T24;
  wire[2:0] T25;
  wire[2:0] T26;
  wire T27;
  wire AcquireTracker_1_io_inner_release_ready;
  wire AcquireTracker_2_io_inner_release_ready;
  wire T28;
  wire T29;
  wire AcquireTracker_3_io_inner_release_ready;
  wire T30;
  wire[1:0] probe_arb_io_out_bits_payload_p_type;
  wire[3:0] probe_arb_io_out_bits_payload_master_xact_id;
  wire[25:0] probe_arb_io_out_bits_payload_addr;
  wire[1:0] probe_arb_io_out_bits_header_dst;
  wire[1:0] probe_arb_io_out_bits_header_src;
  wire probe_arb_io_out_valid;
  wire[3:0] grant_arb_io_out_bits_payload_g_type;
  wire[3:0] grant_arb_io_out_bits_payload_master_xact_id;
  wire[3:0] grant_arb_io_out_bits_payload_client_xact_id;
  wire[511:0] grant_arb_io_out_bits_payload_data;
  wire[1:0] grant_arb_io_out_bits_header_dst;
  wire[1:0] grant_arb_io_out_bits_header_src;
  wire grant_arb_io_out_valid;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;


  assign T0 = io_inner_acquire_valid & T1;
  assign T1 = block_acquires ^ 1'h1;
  assign block_acquires = T2 | AcquireTracker_3_io_has_acquire_conflict;
  assign T2 = T3 | AcquireTracker_2_io_has_acquire_conflict;
  assign T3 = T4 | AcquireTracker_1_io_has_acquire_conflict;
  assign T4 = VoluntaryReleaseTracker_io_has_acquire_conflict | AcquireTracker_0_io_has_acquire_conflict;
  assign T5 = T6;
  assign T6 = {io_incoherent_1, io_incoherent_0};
  assign T7 = io_inner_release_valid & T8;
  assign T8 = release_idx == 4'h4;
  assign release_idx = voluntary ? 4'h0 : io_inner_release_bits_payload_master_xact_id;
  assign voluntary = io_inner_release_bits_payload_r_type == 3'h0;
  assign T9 = T6;
  assign T10 = io_inner_release_valid & T11;
  assign T11 = release_idx == 4'h3;
  assign T12 = T6;
  assign T13 = io_inner_release_valid & T14;
  assign T14 = release_idx == 4'h2;
  assign T15 = T6;
  assign T16 = io_inner_release_valid & T17;
  assign T17 = release_idx == 4'h1;
  assign T18 = T6;
  assign T19 = io_inner_release_valid & T20;
  assign T20 = release_idx == 4'h0;
  assign io_outer_finish_bits_payload_master_xact_id = outer_arb_io_out_finish_bits_payload_master_xact_id;
  assign io_outer_finish_bits_header_dst = outer_arb_io_out_finish_bits_header_dst;
  assign io_outer_finish_bits_header_src = outer_arb_io_out_finish_bits_header_src;
  assign io_outer_finish_valid = outer_arb_io_out_finish_valid;
  assign io_outer_grant_ready = outer_arb_io_out_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = outer_arb_io_out_acquire_bits_payload_atomic_opcode;
  assign io_outer_acquire_bits_payload_subword_addr = outer_arb_io_out_acquire_bits_payload_subword_addr;
  assign io_outer_acquire_bits_payload_write_mask = outer_arb_io_out_acquire_bits_payload_write_mask;
  assign io_outer_acquire_bits_payload_a_type = outer_arb_io_out_acquire_bits_payload_a_type;
  assign io_outer_acquire_bits_payload_data = outer_arb_io_out_acquire_bits_payload_data;
  assign io_outer_acquire_bits_payload_client_xact_id = outer_arb_io_out_acquire_bits_payload_client_xact_id;
  assign io_outer_acquire_bits_payload_addr = outer_arb_io_out_acquire_bits_payload_addr;
  assign io_outer_acquire_bits_header_dst = outer_arb_io_out_acquire_bits_header_dst;
  assign io_outer_acquire_bits_header_src = outer_arb_io_out_acquire_bits_header_src;
  assign io_outer_acquire_valid = outer_arb_io_out_acquire_valid;
  assign io_inner_release_ready = T21;
  assign T21 = T30 ? AcquireTracker_3_io_inner_release_ready : T22;
  assign T22 = T29 ? T27 : T23;
  assign T23 = T24 ? AcquireTracker_0_io_inner_release_ready : VoluntaryReleaseTracker_io_inner_release_ready;
  assign T24 = T25[1'h0:1'h0];
  assign T25 = T26;
  assign T26 = release_idx[2'h2:1'h0];
  assign T27 = T28 ? AcquireTracker_2_io_inner_release_ready : AcquireTracker_1_io_inner_release_ready;
  assign T28 = T25[1'h0:1'h0];
  assign T29 = T25[1'h1:1'h1];
  assign T30 = T25[2'h2:2'h2];
  assign io_inner_probe_bits_payload_p_type = probe_arb_io_out_bits_payload_p_type;
  assign io_inner_probe_bits_payload_master_xact_id = probe_arb_io_out_bits_payload_master_xact_id;
  assign io_inner_probe_bits_payload_addr = probe_arb_io_out_bits_payload_addr;
  assign io_inner_probe_bits_header_dst = probe_arb_io_out_bits_header_dst;
  assign io_inner_probe_bits_header_src = probe_arb_io_out_bits_header_src;
  assign io_inner_probe_valid = probe_arb_io_out_valid;
  assign io_inner_finish_ready = 1'h1;
  assign io_inner_grant_bits_payload_g_type = grant_arb_io_out_bits_payload_g_type;
  assign io_inner_grant_bits_payload_master_xact_id = grant_arb_io_out_bits_payload_master_xact_id;
  assign io_inner_grant_bits_payload_client_xact_id = grant_arb_io_out_bits_payload_client_xact_id;
  assign io_inner_grant_bits_payload_data = grant_arb_io_out_bits_payload_data;
  assign io_inner_grant_bits_header_dst = grant_arb_io_out_bits_header_dst;
  assign io_inner_grant_bits_header_src = grant_arb_io_out_bits_header_src;
  assign io_inner_grant_valid = grant_arb_io_out_valid;
  assign io_inner_acquire_ready = T31;
  assign T31 = T33 & T32;
  assign T32 = block_acquires ^ 1'h1;
  assign T33 = T34 | AcquireTracker_3_io_inner_acquire_ready;
  assign T34 = T35 | AcquireTracker_2_io_inner_acquire_ready;
  assign T35 = T36 | AcquireTracker_1_io_inner_acquire_ready;
  assign T36 = VoluntaryReleaseTracker_io_inner_acquire_ready | AcquireTracker_0_io_inner_acquire_ready;
  VoluntaryReleaseTracker VoluntaryReleaseTracker(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( VoluntaryReleaseTracker_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_0_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_0_ready ),
       .io_inner_grant_valid( VoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( VoluntaryReleaseTracker_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( VoluntaryReleaseTracker_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( VoluntaryReleaseTracker_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_0_ready ),
       .io_inner_probe_valid( VoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_inner_probe_bits_header_src(  )
       //.io_inner_probe_bits_header_dst(  )
       //.io_inner_probe_bits_payload_addr(  )
       //.io_inner_probe_bits_payload_master_xact_id(  )
       //.io_inner_probe_bits_payload_p_type(  )
       .io_inner_release_ready( VoluntaryReleaseTracker_io_inner_release_ready ),
       .io_inner_release_valid( T19 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_outer_acquire_valid( VoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( VoluntaryReleaseTracker_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( VoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_0_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_0_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_0_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_0_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_0_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T18 ),
       .io_has_acquire_conflict( VoluntaryReleaseTracker_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_0 AcquireTracker_0(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_0_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_1_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_1_ready ),
       .io_inner_grant_valid( AcquireTracker_0_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_0_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_0_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_0_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_0_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_1_ready ),
       .io_inner_probe_valid( AcquireTracker_0_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_0_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_0_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_0_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_0_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_0_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_0_io_inner_release_ready ),
       .io_inner_release_valid( T16 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_0_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_0_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_0_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_0_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_0_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_0_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_0_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_0_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_0_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_1_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_1_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_1_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_1_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_1_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T15 ),
       .io_has_acquire_conflict( AcquireTracker_0_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_1 AcquireTracker_1(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_1_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_2_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_2_ready ),
       .io_inner_grant_valid( AcquireTracker_1_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_1_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_1_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_1_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_1_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_2_ready ),
       .io_inner_probe_valid( AcquireTracker_1_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_1_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_1_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_1_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_1_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_1_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_1_io_inner_release_ready ),
       .io_inner_release_valid( T13 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_1_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_1_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_1_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_1_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_1_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_1_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_1_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_1_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_1_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_2_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_2_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_2_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_2_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_2_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_2_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_2_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T12 ),
       .io_has_acquire_conflict( AcquireTracker_1_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_2 AcquireTracker_2(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_2_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_3_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_3_ready ),
       .io_inner_grant_valid( AcquireTracker_2_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_2_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_2_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_2_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_2_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_3_ready ),
       .io_inner_probe_valid( AcquireTracker_2_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_2_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_2_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_2_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_2_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_2_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_2_io_inner_release_ready ),
       .io_inner_release_valid( T10 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_2_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_2_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_2_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_2_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_2_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_2_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_2_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_2_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_2_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_3_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_3_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_3_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_3_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_3_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_3_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_3_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T9 ),
       .io_has_acquire_conflict( AcquireTracker_2_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_3 AcquireTracker_3(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_3_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_4_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_4_ready ),
       .io_inner_grant_valid( AcquireTracker_3_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_3_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_3_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_3_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_3_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_4_ready ),
       .io_inner_probe_valid( AcquireTracker_3_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_3_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_3_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_3_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_3_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_3_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_3_io_inner_release_ready ),
       .io_inner_release_valid( T7 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_3_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_3_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_3_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_3_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_3_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_3_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_3_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_3_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_3_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_4_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_4_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_4_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_4_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_4_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_4_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_4_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T5 ),
       .io_has_acquire_conflict( AcquireTracker_3_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  Arbiter_11 alloc_arb(
       .io_in_4_ready( alloc_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_acquire_ready ),
       //.io_in_4_bits(  )
       .io_in_3_ready( alloc_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_acquire_ready ),
       //.io_in_3_bits(  )
       .io_in_2_ready( alloc_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_acquire_ready ),
       //.io_in_2_bits(  )
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_acquire_ready ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_acquire_ready ),
       //.io_in_0_bits(  )
       .io_out_ready( T0 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign alloc_arb.io_in_4_bits = {1{$random}};
    assign alloc_arb.io_in_3_bits = {1{$random}};
    assign alloc_arb.io_in_2_bits = {1{$random}};
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
  `endif
  Arbiter_12 probe_arb(
       .io_in_4_ready( probe_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_probe_valid ),
       .io_in_4_bits_header_src( AcquireTracker_3_io_inner_probe_bits_header_src ),
       .io_in_4_bits_header_dst( AcquireTracker_3_io_inner_probe_bits_header_dst ),
       .io_in_4_bits_payload_addr( AcquireTracker_3_io_inner_probe_bits_payload_addr ),
       .io_in_4_bits_payload_master_xact_id( AcquireTracker_3_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_4_bits_payload_p_type( AcquireTracker_3_io_inner_probe_bits_payload_p_type ),
       .io_in_3_ready( probe_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_probe_valid ),
       .io_in_3_bits_header_src( AcquireTracker_2_io_inner_probe_bits_header_src ),
       .io_in_3_bits_header_dst( AcquireTracker_2_io_inner_probe_bits_header_dst ),
       .io_in_3_bits_payload_addr( AcquireTracker_2_io_inner_probe_bits_payload_addr ),
       .io_in_3_bits_payload_master_xact_id( AcquireTracker_2_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_3_bits_payload_p_type( AcquireTracker_2_io_inner_probe_bits_payload_p_type ),
       .io_in_2_ready( probe_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_probe_valid ),
       .io_in_2_bits_header_src( AcquireTracker_1_io_inner_probe_bits_header_src ),
       .io_in_2_bits_header_dst( AcquireTracker_1_io_inner_probe_bits_header_dst ),
       .io_in_2_bits_payload_addr( AcquireTracker_1_io_inner_probe_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( AcquireTracker_1_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( AcquireTracker_1_io_inner_probe_bits_payload_p_type ),
       .io_in_1_ready( probe_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_probe_valid ),
       .io_in_1_bits_header_src( AcquireTracker_0_io_inner_probe_bits_header_src ),
       .io_in_1_bits_header_dst( AcquireTracker_0_io_inner_probe_bits_header_dst ),
       .io_in_1_bits_payload_addr( AcquireTracker_0_io_inner_probe_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( AcquireTracker_0_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( AcquireTracker_0_io_inner_probe_bits_payload_p_type ),
       .io_in_0_ready( probe_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_master_xact_id(  )
       //.io_in_0_bits_payload_p_type(  )
       .io_out_ready( io_inner_probe_ready ),
       .io_out_valid( probe_arb_io_out_valid ),
       .io_out_bits_header_src( probe_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( probe_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( probe_arb_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( probe_arb_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( probe_arb_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign probe_arb.io_in_0_bits_header_src = {1{$random}};
    assign probe_arb.io_in_0_bits_header_dst = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_addr = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_master_xact_id = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_p_type = {1{$random}};
  `endif
  Arbiter_13 grant_arb(
       .io_in_4_ready( grant_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_grant_valid ),
       .io_in_4_bits_header_src( AcquireTracker_3_io_inner_grant_bits_header_src ),
       .io_in_4_bits_header_dst( AcquireTracker_3_io_inner_grant_bits_header_dst ),
       .io_in_4_bits_payload_data( AcquireTracker_3_io_inner_grant_bits_payload_data ),
       .io_in_4_bits_payload_client_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_master_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_4_bits_payload_g_type( AcquireTracker_3_io_inner_grant_bits_payload_g_type ),
       .io_in_3_ready( grant_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_grant_valid ),
       .io_in_3_bits_header_src( AcquireTracker_2_io_inner_grant_bits_header_src ),
       .io_in_3_bits_header_dst( AcquireTracker_2_io_inner_grant_bits_header_dst ),
       .io_in_3_bits_payload_data( AcquireTracker_2_io_inner_grant_bits_payload_data ),
       .io_in_3_bits_payload_client_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_master_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_3_bits_payload_g_type( AcquireTracker_2_io_inner_grant_bits_payload_g_type ),
       .io_in_2_ready( grant_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_grant_valid ),
       .io_in_2_bits_header_src( AcquireTracker_1_io_inner_grant_bits_header_src ),
       .io_in_2_bits_header_dst( AcquireTracker_1_io_inner_grant_bits_header_dst ),
       .io_in_2_bits_payload_data( AcquireTracker_1_io_inner_grant_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( AcquireTracker_1_io_inner_grant_bits_payload_g_type ),
       .io_in_1_ready( grant_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_grant_valid ),
       .io_in_1_bits_header_src( AcquireTracker_0_io_inner_grant_bits_header_src ),
       .io_in_1_bits_header_dst( AcquireTracker_0_io_inner_grant_bits_header_dst ),
       .io_in_1_bits_payload_data( AcquireTracker_0_io_inner_grant_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( AcquireTracker_0_io_inner_grant_bits_payload_g_type ),
       .io_in_0_ready( grant_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_in_0_bits_header_src( VoluntaryReleaseTracker_io_inner_grant_bits_header_src ),
       .io_in_0_bits_header_dst( VoluntaryReleaseTracker_io_inner_grant_bits_header_dst ),
       .io_in_0_bits_payload_data( VoluntaryReleaseTracker_io_inner_grant_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type ),
       .io_out_ready( io_inner_grant_ready ),
       .io_out_valid( grant_arb_io_out_valid ),
       .io_out_bits_header_src( grant_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( grant_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_data( grant_arb_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( grant_arb_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( grant_arb_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( grant_arb_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  UncachedTileLinkIOArbiterThatPassesId outer_arb(.clk(clk), .reset(reset),
       .io_in_4_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_in_4_acquire_valid( AcquireTracker_3_io_outer_acquire_valid ),
       .io_in_4_acquire_bits_header_src( AcquireTracker_3_io_outer_acquire_bits_header_src ),
       //.io_in_4_acquire_bits_header_dst(  )
       .io_in_4_acquire_bits_payload_addr( AcquireTracker_3_io_outer_acquire_bits_payload_addr ),
       .io_in_4_acquire_bits_payload_client_xact_id( AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_4_acquire_bits_payload_data( AcquireTracker_3_io_outer_acquire_bits_payload_data ),
       .io_in_4_acquire_bits_payload_a_type( AcquireTracker_3_io_outer_acquire_bits_payload_a_type ),
       .io_in_4_acquire_bits_payload_write_mask( AcquireTracker_3_io_outer_acquire_bits_payload_write_mask ),
       .io_in_4_acquire_bits_payload_subword_addr( AcquireTracker_3_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_4_acquire_bits_payload_atomic_opcode( AcquireTracker_3_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_4_grant_ready( AcquireTracker_3_io_outer_grant_ready ),
       .io_in_4_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_in_4_grant_bits_header_src( outer_arb_io_in_4_grant_bits_header_src ),
       .io_in_4_grant_bits_header_dst( outer_arb_io_in_4_grant_bits_header_dst ),
       .io_in_4_grant_bits_payload_data( outer_arb_io_in_4_grant_bits_payload_data ),
       .io_in_4_grant_bits_payload_client_xact_id( outer_arb_io_in_4_grant_bits_payload_client_xact_id ),
       .io_in_4_grant_bits_payload_master_xact_id( outer_arb_io_in_4_grant_bits_payload_master_xact_id ),
       .io_in_4_grant_bits_payload_g_type( outer_arb_io_in_4_grant_bits_payload_g_type ),
       .io_in_4_finish_ready( outer_arb_io_in_4_finish_ready ),
       //.io_in_4_finish_valid(  )
       //.io_in_4_finish_bits_header_src(  )
       //.io_in_4_finish_bits_header_dst(  )
       //.io_in_4_finish_bits_payload_master_xact_id(  )
       .io_in_3_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_in_3_acquire_valid( AcquireTracker_2_io_outer_acquire_valid ),
       .io_in_3_acquire_bits_header_src( AcquireTracker_2_io_outer_acquire_bits_header_src ),
       //.io_in_3_acquire_bits_header_dst(  )
       .io_in_3_acquire_bits_payload_addr( AcquireTracker_2_io_outer_acquire_bits_payload_addr ),
       .io_in_3_acquire_bits_payload_client_xact_id( AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_3_acquire_bits_payload_data( AcquireTracker_2_io_outer_acquire_bits_payload_data ),
       .io_in_3_acquire_bits_payload_a_type( AcquireTracker_2_io_outer_acquire_bits_payload_a_type ),
       .io_in_3_acquire_bits_payload_write_mask( AcquireTracker_2_io_outer_acquire_bits_payload_write_mask ),
       .io_in_3_acquire_bits_payload_subword_addr( AcquireTracker_2_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_3_acquire_bits_payload_atomic_opcode( AcquireTracker_2_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_3_grant_ready( AcquireTracker_2_io_outer_grant_ready ),
       .io_in_3_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_in_3_grant_bits_header_src( outer_arb_io_in_3_grant_bits_header_src ),
       .io_in_3_grant_bits_header_dst( outer_arb_io_in_3_grant_bits_header_dst ),
       .io_in_3_grant_bits_payload_data( outer_arb_io_in_3_grant_bits_payload_data ),
       .io_in_3_grant_bits_payload_client_xact_id( outer_arb_io_in_3_grant_bits_payload_client_xact_id ),
       .io_in_3_grant_bits_payload_master_xact_id( outer_arb_io_in_3_grant_bits_payload_master_xact_id ),
       .io_in_3_grant_bits_payload_g_type( outer_arb_io_in_3_grant_bits_payload_g_type ),
       .io_in_3_finish_ready( outer_arb_io_in_3_finish_ready ),
       //.io_in_3_finish_valid(  )
       //.io_in_3_finish_bits_header_src(  )
       //.io_in_3_finish_bits_header_dst(  )
       //.io_in_3_finish_bits_payload_master_xact_id(  )
       .io_in_2_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_in_2_acquire_valid( AcquireTracker_1_io_outer_acquire_valid ),
       .io_in_2_acquire_bits_header_src( AcquireTracker_1_io_outer_acquire_bits_header_src ),
       //.io_in_2_acquire_bits_header_dst(  )
       .io_in_2_acquire_bits_payload_addr( AcquireTracker_1_io_outer_acquire_bits_payload_addr ),
       .io_in_2_acquire_bits_payload_client_xact_id( AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_2_acquire_bits_payload_data( AcquireTracker_1_io_outer_acquire_bits_payload_data ),
       .io_in_2_acquire_bits_payload_a_type( AcquireTracker_1_io_outer_acquire_bits_payload_a_type ),
       .io_in_2_acquire_bits_payload_write_mask( AcquireTracker_1_io_outer_acquire_bits_payload_write_mask ),
       .io_in_2_acquire_bits_payload_subword_addr( AcquireTracker_1_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_2_acquire_bits_payload_atomic_opcode( AcquireTracker_1_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_2_grant_ready( AcquireTracker_1_io_outer_grant_ready ),
       .io_in_2_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_in_2_grant_bits_header_src( outer_arb_io_in_2_grant_bits_header_src ),
       .io_in_2_grant_bits_header_dst( outer_arb_io_in_2_grant_bits_header_dst ),
       .io_in_2_grant_bits_payload_data( outer_arb_io_in_2_grant_bits_payload_data ),
       .io_in_2_grant_bits_payload_client_xact_id( outer_arb_io_in_2_grant_bits_payload_client_xact_id ),
       .io_in_2_grant_bits_payload_master_xact_id( outer_arb_io_in_2_grant_bits_payload_master_xact_id ),
       .io_in_2_grant_bits_payload_g_type( outer_arb_io_in_2_grant_bits_payload_g_type ),
       .io_in_2_finish_ready( outer_arb_io_in_2_finish_ready ),
       //.io_in_2_finish_valid(  )
       //.io_in_2_finish_bits_header_src(  )
       //.io_in_2_finish_bits_header_dst(  )
       //.io_in_2_finish_bits_payload_master_xact_id(  )
       .io_in_1_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( AcquireTracker_0_io_outer_acquire_valid ),
       .io_in_1_acquire_bits_header_src( AcquireTracker_0_io_outer_acquire_bits_header_src ),
       //.io_in_1_acquire_bits_header_dst(  )
       .io_in_1_acquire_bits_payload_addr( AcquireTracker_0_io_outer_acquire_bits_payload_addr ),
       .io_in_1_acquire_bits_payload_client_xact_id( AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_1_acquire_bits_payload_data( AcquireTracker_0_io_outer_acquire_bits_payload_data ),
       .io_in_1_acquire_bits_payload_a_type( AcquireTracker_0_io_outer_acquire_bits_payload_a_type ),
       .io_in_1_acquire_bits_payload_write_mask( AcquireTracker_0_io_outer_acquire_bits_payload_write_mask ),
       .io_in_1_acquire_bits_payload_subword_addr( AcquireTracker_0_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_1_acquire_bits_payload_atomic_opcode( AcquireTracker_0_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_1_grant_ready( AcquireTracker_0_io_outer_grant_ready ),
       .io_in_1_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_header_src( outer_arb_io_in_1_grant_bits_header_src ),
       .io_in_1_grant_bits_header_dst( outer_arb_io_in_1_grant_bits_header_dst ),
       .io_in_1_grant_bits_payload_data( outer_arb_io_in_1_grant_bits_payload_data ),
       .io_in_1_grant_bits_payload_client_xact_id( outer_arb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_in_1_grant_bits_payload_master_xact_id( outer_arb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_in_1_grant_bits_payload_g_type( outer_arb_io_in_1_grant_bits_payload_g_type ),
       .io_in_1_finish_ready( outer_arb_io_in_1_finish_ready ),
       //.io_in_1_finish_valid(  )
       //.io_in_1_finish_bits_header_src(  )
       //.io_in_1_finish_bits_header_dst(  )
       //.io_in_1_finish_bits_payload_master_xact_id(  )
       .io_in_0_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( VoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_in_0_acquire_bits_header_src( VoluntaryReleaseTracker_io_outer_acquire_bits_header_src ),
       //.io_in_0_acquire_bits_header_dst(  )
       .io_in_0_acquire_bits_payload_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr ),
       .io_in_0_acquire_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_0_acquire_bits_payload_data( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data ),
       .io_in_0_acquire_bits_payload_a_type( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type ),
       .io_in_0_acquire_bits_payload_write_mask( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_write_mask ),
       .io_in_0_acquire_bits_payload_subword_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_0_acquire_bits_payload_atomic_opcode( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_0_grant_ready( VoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_in_0_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_header_src( outer_arb_io_in_0_grant_bits_header_src ),
       .io_in_0_grant_bits_header_dst( outer_arb_io_in_0_grant_bits_header_dst ),
       .io_in_0_grant_bits_payload_data( outer_arb_io_in_0_grant_bits_payload_data ),
       .io_in_0_grant_bits_payload_client_xact_id( outer_arb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_in_0_grant_bits_payload_master_xact_id( outer_arb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_in_0_grant_bits_payload_g_type( outer_arb_io_in_0_grant_bits_payload_g_type ),
       .io_in_0_finish_ready( outer_arb_io_in_0_finish_ready ),
       //.io_in_0_finish_valid(  )
       //.io_in_0_finish_bits_header_src(  )
       //.io_in_0_finish_bits_header_dst(  )
       //.io_in_0_finish_bits_payload_master_xact_id(  )
       .io_out_acquire_ready( io_outer_acquire_ready ),
       .io_out_acquire_valid( outer_arb_io_out_acquire_valid ),
       .io_out_acquire_bits_header_src( outer_arb_io_out_acquire_bits_header_src ),
       .io_out_acquire_bits_header_dst( outer_arb_io_out_acquire_bits_header_dst ),
       .io_out_acquire_bits_payload_addr( outer_arb_io_out_acquire_bits_payload_addr ),
       .io_out_acquire_bits_payload_client_xact_id( outer_arb_io_out_acquire_bits_payload_client_xact_id ),
       .io_out_acquire_bits_payload_data( outer_arb_io_out_acquire_bits_payload_data ),
       .io_out_acquire_bits_payload_a_type( outer_arb_io_out_acquire_bits_payload_a_type ),
       .io_out_acquire_bits_payload_write_mask( outer_arb_io_out_acquire_bits_payload_write_mask ),
       .io_out_acquire_bits_payload_subword_addr( outer_arb_io_out_acquire_bits_payload_subword_addr ),
       .io_out_acquire_bits_payload_atomic_opcode( outer_arb_io_out_acquire_bits_payload_atomic_opcode ),
       .io_out_grant_ready( outer_arb_io_out_grant_ready ),
       .io_out_grant_valid( io_outer_grant_valid ),
       .io_out_grant_bits_header_src( io_outer_grant_bits_header_src ),
       .io_out_grant_bits_header_dst( io_outer_grant_bits_header_dst ),
       .io_out_grant_bits_payload_data( io_outer_grant_bits_payload_data ),
       .io_out_grant_bits_payload_client_xact_id( io_outer_grant_bits_payload_client_xact_id ),
       .io_out_grant_bits_payload_master_xact_id( io_outer_grant_bits_payload_master_xact_id ),
       .io_out_grant_bits_payload_g_type( io_outer_grant_bits_payload_g_type ),
       .io_out_finish_ready( io_outer_finish_ready ),
       .io_out_finish_valid( outer_arb_io_out_finish_valid ),
       .io_out_finish_bits_header_src( outer_arb_io_out_finish_bits_header_src ),
       .io_out_finish_bits_header_dst( outer_arb_io_out_finish_bits_header_dst ),
       .io_out_finish_bits_payload_master_xact_id( outer_arb_io_out_finish_bits_payload_master_xact_id )
  );
  `ifndef SYNTHESIS
    assign outer_arb.io_in_4_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_4_finish_valid = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_3_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_3_finish_valid = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_2_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_2_finish_valid = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_1_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_1_finish_valid = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_0_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_0_finish_valid = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_payload_master_xact_id = {1{$random}};
  `endif
endmodule

module LockingRRArbiter_0(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [3:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_a_type,
    input [5:0] io_in_2_bits_payload_write_mask,
    input [2:0] io_in_2_bits_payload_subword_addr,
    input [3:0] io_in_2_bits_payload_atomic_opcode,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [3:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [3:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[3:0] io_out_bits_payload_client_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_a_type,
    output[5:0] io_out_bits_payload_write_mask,
    output[2:0] io_out_bits_payload_subword_addr,
    output[3:0] io_out_bits_payload_atomic_opcode,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire T13;
  wire[1:0] T14;
  wire T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire T18;
  wire T19;
  wire[5:0] T20;
  wire[5:0] T21;
  wire T22;
  wire T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  wire T27;
  wire[511:0] T28;
  wire[511:0] T29;
  wire T30;
  wire T31;
  wire[3:0] T32;
  wire[3:0] T33;
  wire T34;
  wire T35;
  wire[25:0] T36;
  wire[25:0] T37;
  wire T38;
  wire T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire ctrl_3;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire ctrl_4;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire ctrl_1;
  wire T72;
  wire T73;
  wire T74;
  wire ctrl_5;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire ctrl_2;
  wire T81;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T9 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T6 = reset ? 2'h0 : T7;
  assign T7 = T8 ? T0 : last_grant;
  assign T8 = io_out_ready & io_out_valid;
  assign T9 = io_in_1_valid & T10;
  assign T10 = last_grant < 2'h1;
  assign io_out_bits_payload_atomic_opcode = T11;
  assign T11 = T15 ? io_in_2_bits_payload_atomic_opcode : T12;
  assign T12 = T13 ? io_in_1_bits_payload_atomic_opcode : io_in_0_bits_payload_atomic_opcode;
  assign T13 = T14[1'h0:1'h0];
  assign T14 = T0;
  assign T15 = T14[1'h1:1'h1];
  assign io_out_bits_payload_subword_addr = T16;
  assign T16 = T19 ? io_in_2_bits_payload_subword_addr : T17;
  assign T17 = T18 ? io_in_1_bits_payload_subword_addr : io_in_0_bits_payload_subword_addr;
  assign T18 = T14[1'h0:1'h0];
  assign T19 = T14[1'h1:1'h1];
  assign io_out_bits_payload_write_mask = T20;
  assign T20 = T23 ? io_in_2_bits_payload_write_mask : T21;
  assign T21 = T22 ? io_in_1_bits_payload_write_mask : io_in_0_bits_payload_write_mask;
  assign T22 = T14[1'h0:1'h0];
  assign T23 = T14[1'h1:1'h1];
  assign io_out_bits_payload_a_type = T24;
  assign T24 = T27 ? io_in_2_bits_payload_a_type : T25;
  assign T25 = T26 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T26 = T14[1'h0:1'h0];
  assign T27 = T14[1'h1:1'h1];
  assign io_out_bits_payload_data = T28;
  assign T28 = T31 ? io_in_2_bits_payload_data : T29;
  assign T29 = T30 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T30 = T14[1'h0:1'h0];
  assign T31 = T14[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T32;
  assign T32 = T35 ? io_in_2_bits_payload_client_xact_id : T33;
  assign T33 = T34 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T34 = T14[1'h0:1'h0];
  assign T35 = T14[1'h1:1'h1];
  assign io_out_bits_payload_addr = T36;
  assign T36 = T39 ? io_in_2_bits_payload_addr : T37;
  assign T37 = T38 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T38 = T14[1'h0:1'h0];
  assign T39 = T14[1'h1:1'h1];
  assign io_out_bits_header_dst = T40;
  assign T40 = T43 ? io_in_2_bits_header_dst : T41;
  assign T41 = T42 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T42 = T14[1'h0:1'h0];
  assign T43 = T14[1'h1:1'h1];
  assign io_out_bits_header_src = T44;
  assign T44 = T47 ? io_in_2_bits_header_src : T45;
  assign T45 = T46 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T46 = T14[1'h0:1'h0];
  assign T47 = T14[1'h1:1'h1];
  assign io_out_valid = T48;
  assign T48 = T51 ? io_in_2_valid : T49;
  assign T49 = T50 ? io_in_1_valid : io_in_0_valid;
  assign T50 = T14[1'h0:1'h0];
  assign T51 = T14[1'h1:1'h1];
  assign io_in_0_ready = T52;
  assign T52 = T53 & io_out_ready;
  assign T53 = T54;
  assign T54 = T63 | ctrl_3;
  assign ctrl_3 = T55 ^ 1'h1;
  assign T55 = T58 | T56;
  assign T56 = io_in_2_valid & T57;
  assign T57 = last_grant < 2'h2;
  assign T58 = T61 | T59;
  assign T59 = io_in_1_valid & T60;
  assign T60 = last_grant < 2'h1;
  assign T61 = io_in_0_valid & T62;
  assign T62 = last_grant < 2'h0;
  assign T63 = last_grant < 2'h0;
  assign io_in_1_ready = T64;
  assign T64 = T65 & io_out_ready;
  assign T65 = T66;
  assign T66 = T70 | ctrl_4;
  assign ctrl_4 = T67 ^ 1'h1;
  assign T67 = T68 | io_in_0_valid;
  assign T68 = T69 | T56;
  assign T69 = T61 | T59;
  assign T70 = ctrl_1 & T71;
  assign T71 = last_grant < 2'h1;
  assign ctrl_1 = T61 ^ 1'h1;
  assign io_in_2_ready = T72;
  assign T72 = T73 & io_out_ready;
  assign T73 = T74;
  assign T74 = T79 | ctrl_5;
  assign ctrl_5 = T75 ^ 1'h1;
  assign T75 = T76 | io_in_1_valid;
  assign T76 = T77 | io_in_0_valid;
  assign T77 = T78 | T56;
  assign T78 = T61 | T59;
  assign T79 = ctrl_2 & T80;
  assign T80 = last_grant < 2'h2;
  assign ctrl_2 = T81 ^ 1'h1;
  assign T81 = T61 | T59;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T8) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_0(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [3:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_a_type,
    input [5:0] io_in_2_bits_payload_write_mask,
    input [2:0] io_in_2_bits_payload_subword_addr,
    input [3:0] io_in_2_bits_payload_atomic_opcode,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [3:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [3:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[3:0] io_out_2_bits_payload_client_xact_id,
    output[511:0] io_out_2_bits_payload_data,
    output[2:0] io_out_2_bits_payload_a_type,
    output[5:0] io_out_2_bits_payload_write_mask,
    output[2:0] io_out_2_bits_payload_subword_addr,
    output[3:0] io_out_2_bits_payload_atomic_opcode,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[3:0] io_out_1_bits_payload_client_xact_id,
    output[511:0] io_out_1_bits_payload_data,
    output[2:0] io_out_1_bits_payload_a_type,
    output[5:0] io_out_1_bits_payload_write_mask,
    output[2:0] io_out_1_bits_payload_subword_addr,
    output[3:0] io_out_1_bits_payload_atomic_opcode,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[3:0] io_out_0_bits_payload_client_xact_id,
    output[511:0] io_out_0_bits_payload_data,
    output[2:0] io_out_0_bits_payload_a_type,
    output[5:0] io_out_0_bits_payload_write_mask,
    output[2:0] io_out_0_bits_payload_subword_addr,
    output[3:0] io_out_0_bits_payload_atomic_opcode
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[3:0] LockingRRArbiter_0_io_out_bits_payload_atomic_opcode;
  wire[2:0] LockingRRArbiter_0_io_out_bits_payload_subword_addr;
  wire[5:0] LockingRRArbiter_0_io_out_bits_payload_write_mask;
  wire[2:0] LockingRRArbiter_0_io_out_bits_payload_a_type;
  wire[511:0] LockingRRArbiter_0_io_out_bits_payload_data;
  wire[3:0] LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[25:0] LockingRRArbiter_0_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_src;
  wire LockingRRArbiter_0_io_out_valid;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_atomic_opcode;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_subword_addr;
  wire[5:0] LockingRRArbiter_1_io_out_bits_payload_write_mask;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_a_type;
  wire[511:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire LockingRRArbiter_1_io_out_valid;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_atomic_opcode;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_subword_addr;
  wire[5:0] LockingRRArbiter_2_io_out_bits_payload_write_mask;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_a_type;
  wire[511:0] LockingRRArbiter_2_io_out_bits_payload_data;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  wire[25:0] LockingRRArbiter_2_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire LockingRRArbiter_2_io_out_valid;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire T26;
  wire T27;
  wire T28;
  wire LockingRRArbiter_0_io_in_0_ready;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire T37;
  wire T38;
  wire T39;
  wire LockingRRArbiter_0_io_in_1_ready;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire T48;
  wire T49;
  wire T50;
  wire LockingRRArbiter_0_io_in_2_ready;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 2'h2;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 2'h2;
  assign T6 = io_in_0_valid & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = io_in_1_valid & T9;
  assign T9 = io_in_1_bits_header_dst == 2'h1;
  assign T10 = io_in_2_valid & T11;
  assign T11 = io_in_2_bits_header_dst == 2'h1;
  assign T12 = io_in_0_valid & T13;
  assign T13 = io_in_0_bits_header_dst == 2'h0;
  assign T14 = io_in_1_valid & T15;
  assign T15 = io_in_1_bits_header_dst == 2'h0;
  assign T16 = io_in_2_valid & T17;
  assign T17 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_atomic_opcode = LockingRRArbiter_0_io_out_bits_payload_atomic_opcode;
  assign io_out_0_bits_payload_subword_addr = LockingRRArbiter_0_io_out_bits_payload_subword_addr;
  assign io_out_0_bits_payload_write_mask = LockingRRArbiter_0_io_out_bits_payload_write_mask;
  assign io_out_0_bits_payload_a_type = LockingRRArbiter_0_io_out_bits_payload_a_type;
  assign io_out_0_bits_payload_data = LockingRRArbiter_0_io_out_bits_payload_data;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_0_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_0_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_0_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_0_io_out_valid;
  assign io_out_1_bits_payload_atomic_opcode = LockingRRArbiter_1_io_out_bits_payload_atomic_opcode;
  assign io_out_1_bits_payload_subword_addr = LockingRRArbiter_1_io_out_bits_payload_subword_addr;
  assign io_out_1_bits_payload_write_mask = LockingRRArbiter_1_io_out_bits_payload_write_mask;
  assign io_out_1_bits_payload_a_type = LockingRRArbiter_1_io_out_bits_payload_a_type;
  assign io_out_1_bits_payload_data = LockingRRArbiter_1_io_out_bits_payload_data;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_1_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_atomic_opcode = LockingRRArbiter_2_io_out_bits_payload_atomic_opcode;
  assign io_out_2_bits_payload_subword_addr = LockingRRArbiter_2_io_out_bits_payload_subword_addr;
  assign io_out_2_bits_payload_write_mask = LockingRRArbiter_2_io_out_bits_payload_write_mask;
  assign io_out_2_bits_payload_a_type = LockingRRArbiter_2_io_out_bits_payload_a_type;
  assign io_out_2_bits_payload_data = LockingRRArbiter_2_io_out_bits_payload_data;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_2_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_in_0_ready = T18;
  assign T18 = T22 | T19;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_2_io_in_0_ready & T21;
  assign T21 = io_in_0_bits_header_dst == 2'h2;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_1_io_in_0_ready & T25;
  assign T25 = io_in_0_bits_header_dst == 2'h1;
  assign T26 = T27;
  assign T27 = LockingRRArbiter_0_io_in_0_ready & T28;
  assign T28 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T29;
  assign T29 = T33 | T30;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_2_io_in_1_ready & T32;
  assign T32 = io_in_1_bits_header_dst == 2'h2;
  assign T33 = T37 | T34;
  assign T34 = T35;
  assign T35 = LockingRRArbiter_1_io_in_1_ready & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h1;
  assign T37 = T38;
  assign T38 = LockingRRArbiter_0_io_in_1_ready & T39;
  assign T39 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T40;
  assign T40 = T44 | T41;
  assign T41 = T42;
  assign T42 = LockingRRArbiter_2_io_in_2_ready & T43;
  assign T43 = io_in_2_bits_header_dst == 2'h2;
  assign T44 = T48 | T45;
  assign T45 = T46;
  assign T46 = LockingRRArbiter_1_io_in_2_ready & T47;
  assign T47 = io_in_2_bits_header_dst == 2'h1;
  assign T48 = T49;
  assign T49 = LockingRRArbiter_0_io_in_2_ready & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_0 LockingRRArbiter_0(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( T16 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_bits_payload_atomic_opcode ),
       .io_in_1_ready( LockingRRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_bits_payload_atomic_opcode ),
       .io_in_0_ready( LockingRRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( T12 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( LockingRRArbiter_0_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( LockingRRArbiter_0_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( LockingRRArbiter_0_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( LockingRRArbiter_0_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  LockingRRArbiter_0 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_bits_payload_atomic_opcode ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T8 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_bits_payload_atomic_opcode ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T6 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_1_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( LockingRRArbiter_1_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( LockingRRArbiter_1_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( LockingRRArbiter_1_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( LockingRRArbiter_1_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  LockingRRArbiter_0 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_bits_payload_atomic_opcode ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_bits_payload_atomic_opcode ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_2_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_2_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( LockingRRArbiter_2_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( LockingRRArbiter_2_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( LockingRRArbiter_2_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( LockingRRArbiter_2_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [3:0] io_in_2_bits_payload_client_xact_id,
    input [3:0] io_in_2_bits_payload_master_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_r_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [3:0] io_in_1_bits_payload_client_xact_id,
    input [3:0] io_in_1_bits_payload_master_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [3:0] io_in_0_bits_payload_client_xact_id,
    input [3:0] io_in_0_bits_payload_master_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[3:0] io_out_bits_payload_client_xact_id,
    output[3:0] io_out_bits_payload_master_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_r_type,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire[1:0] T14;
  wire T15;
  wire[511:0] T16;
  wire[511:0] T17;
  wire T18;
  wire T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T25;
  wire T26;
  wire T27;
  wire[25:0] T28;
  wire[25:0] T29;
  wire T30;
  wire T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire ctrl_3;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire ctrl_4;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire ctrl_1;
  wire T64;
  wire T65;
  wire T66;
  wire ctrl_5;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire ctrl_2;
  wire T73;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T9 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T6 = reset ? 2'h0 : T7;
  assign T7 = T8 ? T0 : last_grant;
  assign T8 = io_out_ready & io_out_valid;
  assign T9 = io_in_1_valid & T10;
  assign T10 = last_grant < 2'h1;
  assign io_out_bits_payload_r_type = T11;
  assign T11 = T15 ? io_in_2_bits_payload_r_type : T12;
  assign T12 = T13 ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign T13 = T14[1'h0:1'h0];
  assign T14 = T0;
  assign T15 = T14[1'h1:1'h1];
  assign io_out_bits_payload_data = T16;
  assign T16 = T19 ? io_in_2_bits_payload_data : T17;
  assign T17 = T18 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T18 = T14[1'h0:1'h0];
  assign T19 = T14[1'h1:1'h1];
  assign io_out_bits_payload_master_xact_id = T20;
  assign T20 = T23 ? io_in_2_bits_payload_master_xact_id : T21;
  assign T21 = T22 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T22 = T14[1'h0:1'h0];
  assign T23 = T14[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T24;
  assign T24 = T27 ? io_in_2_bits_payload_client_xact_id : T25;
  assign T25 = T26 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T26 = T14[1'h0:1'h0];
  assign T27 = T14[1'h1:1'h1];
  assign io_out_bits_payload_addr = T28;
  assign T28 = T31 ? io_in_2_bits_payload_addr : T29;
  assign T29 = T30 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T30 = T14[1'h0:1'h0];
  assign T31 = T14[1'h1:1'h1];
  assign io_out_bits_header_dst = T32;
  assign T32 = T35 ? io_in_2_bits_header_dst : T33;
  assign T33 = T34 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T34 = T14[1'h0:1'h0];
  assign T35 = T14[1'h1:1'h1];
  assign io_out_bits_header_src = T36;
  assign T36 = T39 ? io_in_2_bits_header_src : T37;
  assign T37 = T38 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T38 = T14[1'h0:1'h0];
  assign T39 = T14[1'h1:1'h1];
  assign io_out_valid = T40;
  assign T40 = T43 ? io_in_2_valid : T41;
  assign T41 = T42 ? io_in_1_valid : io_in_0_valid;
  assign T42 = T14[1'h0:1'h0];
  assign T43 = T14[1'h1:1'h1];
  assign io_in_0_ready = T44;
  assign T44 = T45 & io_out_ready;
  assign T45 = T46;
  assign T46 = T55 | ctrl_3;
  assign ctrl_3 = T47 ^ 1'h1;
  assign T47 = T50 | T48;
  assign T48 = io_in_2_valid & T49;
  assign T49 = last_grant < 2'h2;
  assign T50 = T53 | T51;
  assign T51 = io_in_1_valid & T52;
  assign T52 = last_grant < 2'h1;
  assign T53 = io_in_0_valid & T54;
  assign T54 = last_grant < 2'h0;
  assign T55 = last_grant < 2'h0;
  assign io_in_1_ready = T56;
  assign T56 = T57 & io_out_ready;
  assign T57 = T58;
  assign T58 = T62 | ctrl_4;
  assign ctrl_4 = T59 ^ 1'h1;
  assign T59 = T60 | io_in_0_valid;
  assign T60 = T61 | T48;
  assign T61 = T53 | T51;
  assign T62 = ctrl_1 & T63;
  assign T63 = last_grant < 2'h1;
  assign ctrl_1 = T53 ^ 1'h1;
  assign io_in_2_ready = T64;
  assign T64 = T65 & io_out_ready;
  assign T65 = T66;
  assign T66 = T71 | ctrl_5;
  assign ctrl_5 = T67 ^ 1'h1;
  assign T67 = T68 | io_in_1_valid;
  assign T68 = T69 | io_in_0_valid;
  assign T69 = T70 | T48;
  assign T70 = T53 | T51;
  assign T71 = ctrl_2 & T72;
  assign T72 = last_grant < 2'h2;
  assign ctrl_2 = T73 ^ 1'h1;
  assign T73 = T53 | T51;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T8) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [3:0] io_in_2_bits_payload_client_xact_id,
    input [3:0] io_in_2_bits_payload_master_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_r_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [3:0] io_in_1_bits_payload_client_xact_id,
    input [3:0] io_in_1_bits_payload_master_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [3:0] io_in_0_bits_payload_client_xact_id,
    input [3:0] io_in_0_bits_payload_master_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_r_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[3:0] io_out_2_bits_payload_client_xact_id,
    output[3:0] io_out_2_bits_payload_master_xact_id,
    output[511:0] io_out_2_bits_payload_data,
    output[2:0] io_out_2_bits_payload_r_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[3:0] io_out_1_bits_payload_client_xact_id,
    output[3:0] io_out_1_bits_payload_master_xact_id,
    output[511:0] io_out_1_bits_payload_data,
    output[2:0] io_out_1_bits_payload_r_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[3:0] io_out_0_bits_payload_client_xact_id,
    output[3:0] io_out_0_bits_payload_master_xact_id,
    output[511:0] io_out_0_bits_payload_data,
    output[2:0] io_out_0_bits_payload_r_type
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[2:0] LockingRRArbiter_0_io_out_bits_payload_r_type;
  wire[511:0] LockingRRArbiter_0_io_out_bits_payload_data;
  wire[3:0] LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  wire[3:0] LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[25:0] LockingRRArbiter_0_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_src;
  wire LockingRRArbiter_0_io_out_valid;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_r_type;
  wire[511:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire LockingRRArbiter_1_io_out_valid;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_r_type;
  wire[511:0] LockingRRArbiter_2_io_out_bits_payload_data;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  wire[25:0] LockingRRArbiter_2_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire LockingRRArbiter_2_io_out_valid;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire T26;
  wire T27;
  wire T28;
  wire LockingRRArbiter_0_io_in_0_ready;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire T37;
  wire T38;
  wire T39;
  wire LockingRRArbiter_0_io_in_1_ready;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire T48;
  wire T49;
  wire T50;
  wire LockingRRArbiter_0_io_in_2_ready;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 2'h2;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 2'h2;
  assign T6 = io_in_0_valid & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = io_in_1_valid & T9;
  assign T9 = io_in_1_bits_header_dst == 2'h1;
  assign T10 = io_in_2_valid & T11;
  assign T11 = io_in_2_bits_header_dst == 2'h1;
  assign T12 = io_in_0_valid & T13;
  assign T13 = io_in_0_bits_header_dst == 2'h0;
  assign T14 = io_in_1_valid & T15;
  assign T15 = io_in_1_bits_header_dst == 2'h0;
  assign T16 = io_in_2_valid & T17;
  assign T17 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_r_type = LockingRRArbiter_0_io_out_bits_payload_r_type;
  assign io_out_0_bits_payload_data = LockingRRArbiter_0_io_out_bits_payload_data;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_0_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_0_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_0_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_0_io_out_valid;
  assign io_out_1_bits_payload_r_type = LockingRRArbiter_1_io_out_bits_payload_r_type;
  assign io_out_1_bits_payload_data = LockingRRArbiter_1_io_out_bits_payload_data;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_1_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_r_type = LockingRRArbiter_2_io_out_bits_payload_r_type;
  assign io_out_2_bits_payload_data = LockingRRArbiter_2_io_out_bits_payload_data;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_2_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_in_0_ready = T18;
  assign T18 = T22 | T19;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_2_io_in_0_ready & T21;
  assign T21 = io_in_0_bits_header_dst == 2'h2;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_1_io_in_0_ready & T25;
  assign T25 = io_in_0_bits_header_dst == 2'h1;
  assign T26 = T27;
  assign T27 = LockingRRArbiter_0_io_in_0_ready & T28;
  assign T28 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T29;
  assign T29 = T33 | T30;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_2_io_in_1_ready & T32;
  assign T32 = io_in_1_bits_header_dst == 2'h2;
  assign T33 = T37 | T34;
  assign T34 = T35;
  assign T35 = LockingRRArbiter_1_io_in_1_ready & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h1;
  assign T37 = T38;
  assign T38 = LockingRRArbiter_0_io_in_1_ready & T39;
  assign T39 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T40;
  assign T40 = T44 | T41;
  assign T41 = T42;
  assign T42 = LockingRRArbiter_2_io_in_2_ready & T43;
  assign T43 = io_in_2_bits_header_dst == 2'h2;
  assign T44 = T48 | T45;
  assign T45 = T46;
  assign T46 = LockingRRArbiter_1_io_in_2_ready & T47;
  assign T47 = io_in_2_bits_header_dst == 2'h1;
  assign T48 = T49;
  assign T49 = LockingRRArbiter_0_io_in_2_ready & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_1 LockingRRArbiter_0(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( T16 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( T12 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_0_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_0_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_1 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T8 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T6 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_1_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_1_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_1_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_1 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_2_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_2_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_2_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_2_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_2(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [3:0] io_in_2_bits_payload_master_xact_id,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [3:0] io_in_1_bits_payload_master_xact_id,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [3:0] io_in_0_bits_payload_master_xact_id,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[3:0] io_out_bits_payload_master_xact_id,
    output[1:0] io_out_bits_payload_p_type,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire[1:0] T14;
  wire T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire T18;
  wire T19;
  wire[25:0] T20;
  wire[25:0] T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire ctrl_3;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire ctrl_4;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire ctrl_1;
  wire T56;
  wire T57;
  wire T58;
  wire ctrl_5;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire ctrl_2;
  wire T65;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T9 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T6 = reset ? 2'h0 : T7;
  assign T7 = T8 ? T0 : last_grant;
  assign T8 = io_out_ready & io_out_valid;
  assign T9 = io_in_1_valid & T10;
  assign T10 = last_grant < 2'h1;
  assign io_out_bits_payload_p_type = T11;
  assign T11 = T15 ? io_in_2_bits_payload_p_type : T12;
  assign T12 = T13 ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign T13 = T14[1'h0:1'h0];
  assign T14 = T0;
  assign T15 = T14[1'h1:1'h1];
  assign io_out_bits_payload_master_xact_id = T16;
  assign T16 = T19 ? io_in_2_bits_payload_master_xact_id : T17;
  assign T17 = T18 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T18 = T14[1'h0:1'h0];
  assign T19 = T14[1'h1:1'h1];
  assign io_out_bits_payload_addr = T20;
  assign T20 = T23 ? io_in_2_bits_payload_addr : T21;
  assign T21 = T22 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T22 = T14[1'h0:1'h0];
  assign T23 = T14[1'h1:1'h1];
  assign io_out_bits_header_dst = T24;
  assign T24 = T27 ? io_in_2_bits_header_dst : T25;
  assign T25 = T26 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T26 = T14[1'h0:1'h0];
  assign T27 = T14[1'h1:1'h1];
  assign io_out_bits_header_src = T28;
  assign T28 = T31 ? io_in_2_bits_header_src : T29;
  assign T29 = T30 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T30 = T14[1'h0:1'h0];
  assign T31 = T14[1'h1:1'h1];
  assign io_out_valid = T32;
  assign T32 = T35 ? io_in_2_valid : T33;
  assign T33 = T34 ? io_in_1_valid : io_in_0_valid;
  assign T34 = T14[1'h0:1'h0];
  assign T35 = T14[1'h1:1'h1];
  assign io_in_0_ready = T36;
  assign T36 = T37 & io_out_ready;
  assign T37 = T38;
  assign T38 = T47 | ctrl_3;
  assign ctrl_3 = T39 ^ 1'h1;
  assign T39 = T42 | T40;
  assign T40 = io_in_2_valid & T41;
  assign T41 = last_grant < 2'h2;
  assign T42 = T45 | T43;
  assign T43 = io_in_1_valid & T44;
  assign T44 = last_grant < 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = last_grant < 2'h0;
  assign T47 = last_grant < 2'h0;
  assign io_in_1_ready = T48;
  assign T48 = T49 & io_out_ready;
  assign T49 = T50;
  assign T50 = T54 | ctrl_4;
  assign ctrl_4 = T51 ^ 1'h1;
  assign T51 = T52 | io_in_0_valid;
  assign T52 = T53 | T40;
  assign T53 = T45 | T43;
  assign T54 = ctrl_1 & T55;
  assign T55 = last_grant < 2'h1;
  assign ctrl_1 = T45 ^ 1'h1;
  assign io_in_2_ready = T56;
  assign T56 = T57 & io_out_ready;
  assign T57 = T58;
  assign T58 = T63 | ctrl_5;
  assign ctrl_5 = T59 ^ 1'h1;
  assign T59 = T60 | io_in_1_valid;
  assign T60 = T61 | io_in_0_valid;
  assign T61 = T62 | T40;
  assign T62 = T45 | T43;
  assign T63 = ctrl_2 & T64;
  assign T64 = last_grant < 2'h2;
  assign ctrl_2 = T65 ^ 1'h1;
  assign T65 = T45 | T43;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T8) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_2(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [3:0] io_in_2_bits_payload_master_xact_id,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [3:0] io_in_1_bits_payload_master_xact_id,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [3:0] io_in_0_bits_payload_master_xact_id,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[3:0] io_out_2_bits_payload_master_xact_id,
    output[1:0] io_out_2_bits_payload_p_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[3:0] io_out_1_bits_payload_master_xact_id,
    output[1:0] io_out_1_bits_payload_p_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[3:0] io_out_0_bits_payload_master_xact_id,
    output[1:0] io_out_0_bits_payload_p_type
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[1:0] LockingRRArbiter_0_io_out_bits_payload_p_type;
  wire[3:0] LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  wire[25:0] LockingRRArbiter_0_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_src;
  wire LockingRRArbiter_0_io_out_valid;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_p_type;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire LockingRRArbiter_1_io_out_valid;
  wire[1:0] LockingRRArbiter_2_io_out_bits_payload_p_type;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  wire[25:0] LockingRRArbiter_2_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire LockingRRArbiter_2_io_out_valid;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire T26;
  wire T27;
  wire T28;
  wire LockingRRArbiter_0_io_in_0_ready;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire T37;
  wire T38;
  wire T39;
  wire LockingRRArbiter_0_io_in_1_ready;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire T48;
  wire T49;
  wire T50;
  wire LockingRRArbiter_0_io_in_2_ready;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 2'h2;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 2'h2;
  assign T6 = io_in_0_valid & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = io_in_1_valid & T9;
  assign T9 = io_in_1_bits_header_dst == 2'h1;
  assign T10 = io_in_2_valid & T11;
  assign T11 = io_in_2_bits_header_dst == 2'h1;
  assign T12 = io_in_0_valid & T13;
  assign T13 = io_in_0_bits_header_dst == 2'h0;
  assign T14 = io_in_1_valid & T15;
  assign T15 = io_in_1_bits_header_dst == 2'h0;
  assign T16 = io_in_2_valid & T17;
  assign T17 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_p_type = LockingRRArbiter_0_io_out_bits_payload_p_type;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_0_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_0_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_0_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_0_io_out_valid;
  assign io_out_1_bits_payload_p_type = LockingRRArbiter_1_io_out_bits_payload_p_type;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_1_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_p_type = LockingRRArbiter_2_io_out_bits_payload_p_type;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_2_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_in_0_ready = T18;
  assign T18 = T22 | T19;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_2_io_in_0_ready & T21;
  assign T21 = io_in_0_bits_header_dst == 2'h2;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_1_io_in_0_ready & T25;
  assign T25 = io_in_0_bits_header_dst == 2'h1;
  assign T26 = T27;
  assign T27 = LockingRRArbiter_0_io_in_0_ready & T28;
  assign T28 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T29;
  assign T29 = T33 | T30;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_2_io_in_1_ready & T32;
  assign T32 = io_in_1_bits_header_dst == 2'h2;
  assign T33 = T37 | T34;
  assign T34 = T35;
  assign T35 = LockingRRArbiter_1_io_in_1_ready & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h1;
  assign T37 = T38;
  assign T38 = LockingRRArbiter_0_io_in_1_ready & T39;
  assign T39 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T40;
  assign T40 = T44 | T41;
  assign T41 = T42;
  assign T42 = LockingRRArbiter_2_io_in_2_ready & T43;
  assign T43 = io_in_2_bits_header_dst == 2'h2;
  assign T44 = T48 | T45;
  assign T45 = T46;
  assign T46 = LockingRRArbiter_1_io_in_2_ready & T47;
  assign T47 = io_in_2_bits_header_dst == 2'h1;
  assign T48 = T49;
  assign T49 = LockingRRArbiter_0_io_in_2_ready & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_2 LockingRRArbiter_0(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( T16 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( T12 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_0_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( LockingRRArbiter_0_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_2 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T8 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T6 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_1_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_1_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( LockingRRArbiter_1_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_2 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_2_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_2_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( LockingRRArbiter_2_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_3(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [511:0] io_in_2_bits_payload_data,
    input [3:0] io_in_2_bits_payload_client_xact_id,
    input [3:0] io_in_2_bits_payload_master_xact_id,
    input [3:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [511:0] io_in_1_bits_payload_data,
    input [3:0] io_in_1_bits_payload_client_xact_id,
    input [3:0] io_in_1_bits_payload_master_xact_id,
    input [3:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [511:0] io_in_0_bits_payload_data,
    input [3:0] io_in_0_bits_payload_client_xact_id,
    input [3:0] io_in_0_bits_payload_master_xact_id,
    input [3:0] io_in_0_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[3:0] io_out_bits_payload_client_xact_id,
    output[3:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire T13;
  wire[1:0] T14;
  wire T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire T18;
  wire T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire T22;
  wire T23;
  wire[511:0] T24;
  wire[511:0] T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire ctrl_3;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire ctrl_4;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire ctrl_1;
  wire T60;
  wire T61;
  wire T62;
  wire ctrl_5;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire ctrl_2;
  wire T69;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T9 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T6 = reset ? 2'h0 : T7;
  assign T7 = T8 ? T0 : last_grant;
  assign T8 = io_out_ready & io_out_valid;
  assign T9 = io_in_1_valid & T10;
  assign T10 = last_grant < 2'h1;
  assign io_out_bits_payload_g_type = T11;
  assign T11 = T15 ? io_in_2_bits_payload_g_type : T12;
  assign T12 = T13 ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign T13 = T14[1'h0:1'h0];
  assign T14 = T0;
  assign T15 = T14[1'h1:1'h1];
  assign io_out_bits_payload_master_xact_id = T16;
  assign T16 = T19 ? io_in_2_bits_payload_master_xact_id : T17;
  assign T17 = T18 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T18 = T14[1'h0:1'h0];
  assign T19 = T14[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T20;
  assign T20 = T23 ? io_in_2_bits_payload_client_xact_id : T21;
  assign T21 = T22 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T22 = T14[1'h0:1'h0];
  assign T23 = T14[1'h1:1'h1];
  assign io_out_bits_payload_data = T24;
  assign T24 = T27 ? io_in_2_bits_payload_data : T25;
  assign T25 = T26 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T26 = T14[1'h0:1'h0];
  assign T27 = T14[1'h1:1'h1];
  assign io_out_bits_header_dst = T28;
  assign T28 = T31 ? io_in_2_bits_header_dst : T29;
  assign T29 = T30 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T30 = T14[1'h0:1'h0];
  assign T31 = T14[1'h1:1'h1];
  assign io_out_bits_header_src = T32;
  assign T32 = T35 ? io_in_2_bits_header_src : T33;
  assign T33 = T34 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T34 = T14[1'h0:1'h0];
  assign T35 = T14[1'h1:1'h1];
  assign io_out_valid = T36;
  assign T36 = T39 ? io_in_2_valid : T37;
  assign T37 = T38 ? io_in_1_valid : io_in_0_valid;
  assign T38 = T14[1'h0:1'h0];
  assign T39 = T14[1'h1:1'h1];
  assign io_in_0_ready = T40;
  assign T40 = T41 & io_out_ready;
  assign T41 = T42;
  assign T42 = T51 | ctrl_3;
  assign ctrl_3 = T43 ^ 1'h1;
  assign T43 = T46 | T44;
  assign T44 = io_in_2_valid & T45;
  assign T45 = last_grant < 2'h2;
  assign T46 = T49 | T47;
  assign T47 = io_in_1_valid & T48;
  assign T48 = last_grant < 2'h1;
  assign T49 = io_in_0_valid & T50;
  assign T50 = last_grant < 2'h0;
  assign T51 = last_grant < 2'h0;
  assign io_in_1_ready = T52;
  assign T52 = T53 & io_out_ready;
  assign T53 = T54;
  assign T54 = T58 | ctrl_4;
  assign ctrl_4 = T55 ^ 1'h1;
  assign T55 = T56 | io_in_0_valid;
  assign T56 = T57 | T44;
  assign T57 = T49 | T47;
  assign T58 = ctrl_1 & T59;
  assign T59 = last_grant < 2'h1;
  assign ctrl_1 = T49 ^ 1'h1;
  assign io_in_2_ready = T60;
  assign T60 = T61 & io_out_ready;
  assign T61 = T62;
  assign T62 = T67 | ctrl_5;
  assign ctrl_5 = T63 ^ 1'h1;
  assign T63 = T64 | io_in_1_valid;
  assign T64 = T65 | io_in_0_valid;
  assign T65 = T66 | T44;
  assign T66 = T49 | T47;
  assign T67 = ctrl_2 & T68;
  assign T68 = last_grant < 2'h2;
  assign ctrl_2 = T69 ^ 1'h1;
  assign T69 = T49 | T47;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T8) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_3(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [511:0] io_in_2_bits_payload_data,
    input [3:0] io_in_2_bits_payload_client_xact_id,
    input [3:0] io_in_2_bits_payload_master_xact_id,
    input [3:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [511:0] io_in_1_bits_payload_data,
    input [3:0] io_in_1_bits_payload_client_xact_id,
    input [3:0] io_in_1_bits_payload_master_xact_id,
    input [3:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [511:0] io_in_0_bits_payload_data,
    input [3:0] io_in_0_bits_payload_client_xact_id,
    input [3:0] io_in_0_bits_payload_master_xact_id,
    input [3:0] io_in_0_bits_payload_g_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[511:0] io_out_2_bits_payload_data,
    output[3:0] io_out_2_bits_payload_client_xact_id,
    output[3:0] io_out_2_bits_payload_master_xact_id,
    output[3:0] io_out_2_bits_payload_g_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[511:0] io_out_1_bits_payload_data,
    output[3:0] io_out_1_bits_payload_client_xact_id,
    output[3:0] io_out_1_bits_payload_master_xact_id,
    output[3:0] io_out_1_bits_payload_g_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[511:0] io_out_0_bits_payload_data,
    output[3:0] io_out_0_bits_payload_client_xact_id,
    output[3:0] io_out_0_bits_payload_master_xact_id,
    output[3:0] io_out_0_bits_payload_g_type
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[3:0] LockingRRArbiter_0_io_out_bits_payload_g_type;
  wire[3:0] LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  wire[3:0] LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_0_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_src;
  wire LockingRRArbiter_0_io_out_valid;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_g_type;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire LockingRRArbiter_1_io_out_valid;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_g_type;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_2_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire LockingRRArbiter_2_io_out_valid;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire T26;
  wire T27;
  wire T28;
  wire LockingRRArbiter_0_io_in_0_ready;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire T37;
  wire T38;
  wire T39;
  wire LockingRRArbiter_0_io_in_1_ready;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire T48;
  wire T49;
  wire T50;
  wire LockingRRArbiter_0_io_in_2_ready;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 2'h2;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 2'h2;
  assign T6 = io_in_0_valid & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = io_in_1_valid & T9;
  assign T9 = io_in_1_bits_header_dst == 2'h1;
  assign T10 = io_in_2_valid & T11;
  assign T11 = io_in_2_bits_header_dst == 2'h1;
  assign T12 = io_in_0_valid & T13;
  assign T13 = io_in_0_bits_header_dst == 2'h0;
  assign T14 = io_in_1_valid & T15;
  assign T15 = io_in_1_bits_header_dst == 2'h0;
  assign T16 = io_in_2_valid & T17;
  assign T17 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_g_type = LockingRRArbiter_0_io_out_bits_payload_g_type;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_data = LockingRRArbiter_0_io_out_bits_payload_data;
  assign io_out_0_bits_header_dst = LockingRRArbiter_0_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_0_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_0_io_out_valid;
  assign io_out_1_bits_payload_g_type = LockingRRArbiter_1_io_out_bits_payload_g_type;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_data = LockingRRArbiter_1_io_out_bits_payload_data;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_g_type = LockingRRArbiter_2_io_out_bits_payload_g_type;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_data = LockingRRArbiter_2_io_out_bits_payload_data;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_in_0_ready = T18;
  assign T18 = T22 | T19;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_2_io_in_0_ready & T21;
  assign T21 = io_in_0_bits_header_dst == 2'h2;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_1_io_in_0_ready & T25;
  assign T25 = io_in_0_bits_header_dst == 2'h1;
  assign T26 = T27;
  assign T27 = LockingRRArbiter_0_io_in_0_ready & T28;
  assign T28 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T29;
  assign T29 = T33 | T30;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_2_io_in_1_ready & T32;
  assign T32 = io_in_1_bits_header_dst == 2'h2;
  assign T33 = T37 | T34;
  assign T34 = T35;
  assign T35 = LockingRRArbiter_1_io_in_1_ready & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h1;
  assign T37 = T38;
  assign T38 = LockingRRArbiter_0_io_in_1_ready & T39;
  assign T39 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T40;
  assign T40 = T44 | T41;
  assign T41 = T42;
  assign T42 = LockingRRArbiter_2_io_in_2_ready & T43;
  assign T43 = io_in_2_bits_header_dst == 2'h2;
  assign T44 = T48 | T45;
  assign T45 = T46;
  assign T46 = LockingRRArbiter_1_io_in_2_ready & T47;
  assign T47 = io_in_2_bits_header_dst == 2'h1;
  assign T48 = T49;
  assign T49 = LockingRRArbiter_0_io_in_2_ready & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_3 LockingRRArbiter_0(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( T16 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( T12 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_0_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( LockingRRArbiter_0_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_3 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T8 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T6 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_1_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( LockingRRArbiter_1_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_3 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_2_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_2_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( LockingRRArbiter_2_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_4(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [3:0] io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [3:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [3:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[3:0] io_out_bits_payload_master_xact_id,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire T13;
  wire[1:0] T14;
  wire T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire ctrl_3;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire ctrl_4;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire ctrl_1;
  wire T48;
  wire T49;
  wire T50;
  wire ctrl_5;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire ctrl_2;
  wire T57;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T9 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T6 = reset ? 2'h0 : T7;
  assign T7 = T8 ? T0 : last_grant;
  assign T8 = io_out_ready & io_out_valid;
  assign T9 = io_in_1_valid & T10;
  assign T10 = last_grant < 2'h1;
  assign io_out_bits_payload_master_xact_id = T11;
  assign T11 = T15 ? io_in_2_bits_payload_master_xact_id : T12;
  assign T12 = T13 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T13 = T14[1'h0:1'h0];
  assign T14 = T0;
  assign T15 = T14[1'h1:1'h1];
  assign io_out_bits_header_dst = T16;
  assign T16 = T19 ? io_in_2_bits_header_dst : T17;
  assign T17 = T18 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T18 = T14[1'h0:1'h0];
  assign T19 = T14[1'h1:1'h1];
  assign io_out_bits_header_src = T20;
  assign T20 = T23 ? io_in_2_bits_header_src : T21;
  assign T21 = T22 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T22 = T14[1'h0:1'h0];
  assign T23 = T14[1'h1:1'h1];
  assign io_out_valid = T24;
  assign T24 = T27 ? io_in_2_valid : T25;
  assign T25 = T26 ? io_in_1_valid : io_in_0_valid;
  assign T26 = T14[1'h0:1'h0];
  assign T27 = T14[1'h1:1'h1];
  assign io_in_0_ready = T28;
  assign T28 = T29 & io_out_ready;
  assign T29 = T30;
  assign T30 = T39 | ctrl_3;
  assign ctrl_3 = T31 ^ 1'h1;
  assign T31 = T34 | T32;
  assign T32 = io_in_2_valid & T33;
  assign T33 = last_grant < 2'h2;
  assign T34 = T37 | T35;
  assign T35 = io_in_1_valid & T36;
  assign T36 = last_grant < 2'h1;
  assign T37 = io_in_0_valid & T38;
  assign T38 = last_grant < 2'h0;
  assign T39 = last_grant < 2'h0;
  assign io_in_1_ready = T40;
  assign T40 = T41 & io_out_ready;
  assign T41 = T42;
  assign T42 = T46 | ctrl_4;
  assign ctrl_4 = T43 ^ 1'h1;
  assign T43 = T44 | io_in_0_valid;
  assign T44 = T45 | T32;
  assign T45 = T37 | T35;
  assign T46 = ctrl_1 & T47;
  assign T47 = last_grant < 2'h1;
  assign ctrl_1 = T37 ^ 1'h1;
  assign io_in_2_ready = T48;
  assign T48 = T49 & io_out_ready;
  assign T49 = T50;
  assign T50 = T55 | ctrl_5;
  assign ctrl_5 = T51 ^ 1'h1;
  assign T51 = T52 | io_in_1_valid;
  assign T52 = T53 | io_in_0_valid;
  assign T53 = T54 | T32;
  assign T54 = T37 | T35;
  assign T55 = ctrl_2 & T56;
  assign T56 = last_grant < 2'h2;
  assign ctrl_2 = T57 ^ 1'h1;
  assign T57 = T37 | T35;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T8) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_4(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [3:0] io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [3:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [3:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[3:0] io_out_2_bits_payload_master_xact_id,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[3:0] io_out_1_bits_payload_master_xact_id,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[3:0] io_out_0_bits_payload_master_xact_id
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[3:0] LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_src;
  wire LockingRRArbiter_0_io_out_valid;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire LockingRRArbiter_1_io_out_valid;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire LockingRRArbiter_2_io_out_valid;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire T26;
  wire T27;
  wire T28;
  wire LockingRRArbiter_0_io_in_0_ready;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire T37;
  wire T38;
  wire T39;
  wire LockingRRArbiter_0_io_in_1_ready;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire T48;
  wire T49;
  wire T50;
  wire LockingRRArbiter_0_io_in_2_ready;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 2'h2;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 2'h2;
  assign T6 = io_in_0_valid & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = io_in_1_valid & T9;
  assign T9 = io_in_1_bits_header_dst == 2'h1;
  assign T10 = io_in_2_valid & T11;
  assign T11 = io_in_2_bits_header_dst == 2'h1;
  assign T12 = io_in_0_valid & T13;
  assign T13 = io_in_0_bits_header_dst == 2'h0;
  assign T14 = io_in_1_valid & T15;
  assign T15 = io_in_1_bits_header_dst == 2'h0;
  assign T16 = io_in_2_valid & T17;
  assign T17 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_header_dst = LockingRRArbiter_0_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_0_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_0_io_out_valid;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_in_0_ready = T18;
  assign T18 = T22 | T19;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_2_io_in_0_ready & T21;
  assign T21 = io_in_0_bits_header_dst == 2'h2;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_1_io_in_0_ready & T25;
  assign T25 = io_in_0_bits_header_dst == 2'h1;
  assign T26 = T27;
  assign T27 = LockingRRArbiter_0_io_in_0_ready & T28;
  assign T28 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T29;
  assign T29 = T33 | T30;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_2_io_in_1_ready & T32;
  assign T32 = io_in_1_bits_header_dst == 2'h2;
  assign T33 = T37 | T34;
  assign T34 = T35;
  assign T35 = LockingRRArbiter_1_io_in_1_ready & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h1;
  assign T37 = T38;
  assign T38 = LockingRRArbiter_0_io_in_1_ready & T39;
  assign T39 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T40;
  assign T40 = T44 | T41;
  assign T41 = T42;
  assign T42 = LockingRRArbiter_2_io_in_2_ready & T43;
  assign T43 = io_in_2_bits_header_dst == 2'h2;
  assign T44 = T48 | T45;
  assign T45 = T46;
  assign T46 = LockingRRArbiter_1_io_in_2_ready & T47;
  assign T47 = io_in_2_bits_header_dst == 2'h1;
  assign T48 = T49;
  assign T49 = LockingRRArbiter_0_io_in_2_ready & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_4 LockingRRArbiter_0(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( T16 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_1_ready( LockingRRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_0_ready( LockingRRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( T12 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_0_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_4 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T8 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T6 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_1_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_4 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_2_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
endmodule

module ReferenceChipCrossbarNetwork(input clk, input reset,
    output io_clients_1_acquire_ready,
    input  io_clients_1_acquire_valid,
    input [1:0] io_clients_1_acquire_bits_header_src,
    input [1:0] io_clients_1_acquire_bits_header_dst,
    input [25:0] io_clients_1_acquire_bits_payload_addr,
    input [3:0] io_clients_1_acquire_bits_payload_client_xact_id,
    input [511:0] io_clients_1_acquire_bits_payload_data,
    input [2:0] io_clients_1_acquire_bits_payload_a_type,
    input [5:0] io_clients_1_acquire_bits_payload_write_mask,
    input [2:0] io_clients_1_acquire_bits_payload_subword_addr,
    input [3:0] io_clients_1_acquire_bits_payload_atomic_opcode,
    input  io_clients_1_grant_ready,
    output io_clients_1_grant_valid,
    output[1:0] io_clients_1_grant_bits_header_src,
    output[1:0] io_clients_1_grant_bits_header_dst,
    output[511:0] io_clients_1_grant_bits_payload_data,
    output[3:0] io_clients_1_grant_bits_payload_client_xact_id,
    output[3:0] io_clients_1_grant_bits_payload_master_xact_id,
    output[3:0] io_clients_1_grant_bits_payload_g_type,
    output io_clients_1_finish_ready,
    input  io_clients_1_finish_valid,
    input [1:0] io_clients_1_finish_bits_header_src,
    input [1:0] io_clients_1_finish_bits_header_dst,
    input [3:0] io_clients_1_finish_bits_payload_master_xact_id,
    input  io_clients_1_probe_ready,
    output io_clients_1_probe_valid,
    output[1:0] io_clients_1_probe_bits_header_src,
    output[1:0] io_clients_1_probe_bits_header_dst,
    output[25:0] io_clients_1_probe_bits_payload_addr,
    output[3:0] io_clients_1_probe_bits_payload_master_xact_id,
    output[1:0] io_clients_1_probe_bits_payload_p_type,
    output io_clients_1_release_ready,
    input  io_clients_1_release_valid,
    input [1:0] io_clients_1_release_bits_header_src,
    input [1:0] io_clients_1_release_bits_header_dst,
    input [25:0] io_clients_1_release_bits_payload_addr,
    input [3:0] io_clients_1_release_bits_payload_client_xact_id,
    input [3:0] io_clients_1_release_bits_payload_master_xact_id,
    input [511:0] io_clients_1_release_bits_payload_data,
    input [2:0] io_clients_1_release_bits_payload_r_type,
    output io_clients_0_acquire_ready,
    input  io_clients_0_acquire_valid,
    input [1:0] io_clients_0_acquire_bits_header_src,
    input [1:0] io_clients_0_acquire_bits_header_dst,
    input [25:0] io_clients_0_acquire_bits_payload_addr,
    input [3:0] io_clients_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_clients_0_acquire_bits_payload_data,
    input [2:0] io_clients_0_acquire_bits_payload_a_type,
    input [5:0] io_clients_0_acquire_bits_payload_write_mask,
    input [2:0] io_clients_0_acquire_bits_payload_subword_addr,
    input [3:0] io_clients_0_acquire_bits_payload_atomic_opcode,
    input  io_clients_0_grant_ready,
    output io_clients_0_grant_valid,
    output[1:0] io_clients_0_grant_bits_header_src,
    output[1:0] io_clients_0_grant_bits_header_dst,
    output[511:0] io_clients_0_grant_bits_payload_data,
    output[3:0] io_clients_0_grant_bits_payload_client_xact_id,
    output[3:0] io_clients_0_grant_bits_payload_master_xact_id,
    output[3:0] io_clients_0_grant_bits_payload_g_type,
    output io_clients_0_finish_ready,
    input  io_clients_0_finish_valid,
    input [1:0] io_clients_0_finish_bits_header_src,
    input [1:0] io_clients_0_finish_bits_header_dst,
    input [3:0] io_clients_0_finish_bits_payload_master_xact_id,
    input  io_clients_0_probe_ready,
    output io_clients_0_probe_valid,
    output[1:0] io_clients_0_probe_bits_header_src,
    output[1:0] io_clients_0_probe_bits_header_dst,
    output[25:0] io_clients_0_probe_bits_payload_addr,
    output[3:0] io_clients_0_probe_bits_payload_master_xact_id,
    output[1:0] io_clients_0_probe_bits_payload_p_type,
    output io_clients_0_release_ready,
    input  io_clients_0_release_valid,
    input [1:0] io_clients_0_release_bits_header_src,
    input [1:0] io_clients_0_release_bits_header_dst,
    input [25:0] io_clients_0_release_bits_payload_addr,
    input [3:0] io_clients_0_release_bits_payload_client_xact_id,
    input [3:0] io_clients_0_release_bits_payload_master_xact_id,
    input [511:0] io_clients_0_release_bits_payload_data,
    input [2:0] io_clients_0_release_bits_payload_r_type,
    input  io_masters_0_acquire_ready,
    output io_masters_0_acquire_valid,
    output[1:0] io_masters_0_acquire_bits_header_src,
    output[1:0] io_masters_0_acquire_bits_header_dst,
    output[25:0] io_masters_0_acquire_bits_payload_addr,
    output[3:0] io_masters_0_acquire_bits_payload_client_xact_id,
    output[511:0] io_masters_0_acquire_bits_payload_data,
    output[2:0] io_masters_0_acquire_bits_payload_a_type,
    output[5:0] io_masters_0_acquire_bits_payload_write_mask,
    output[2:0] io_masters_0_acquire_bits_payload_subword_addr,
    output[3:0] io_masters_0_acquire_bits_payload_atomic_opcode,
    output io_masters_0_grant_ready,
    input  io_masters_0_grant_valid,
    input [1:0] io_masters_0_grant_bits_header_src,
    input [1:0] io_masters_0_grant_bits_header_dst,
    input [511:0] io_masters_0_grant_bits_payload_data,
    input [3:0] io_masters_0_grant_bits_payload_client_xact_id,
    input [3:0] io_masters_0_grant_bits_payload_master_xact_id,
    input [3:0] io_masters_0_grant_bits_payload_g_type,
    input  io_masters_0_finish_ready,
    output io_masters_0_finish_valid,
    output[1:0] io_masters_0_finish_bits_header_src,
    output[1:0] io_masters_0_finish_bits_header_dst,
    output[3:0] io_masters_0_finish_bits_payload_master_xact_id,
    output io_masters_0_probe_ready,
    input  io_masters_0_probe_valid,
    input [1:0] io_masters_0_probe_bits_header_src,
    input [1:0] io_masters_0_probe_bits_header_dst,
    input [25:0] io_masters_0_probe_bits_payload_addr,
    input [3:0] io_masters_0_probe_bits_payload_master_xact_id,
    input [1:0] io_masters_0_probe_bits_payload_p_type,
    input  io_masters_0_release_ready,
    output io_masters_0_release_valid,
    output[1:0] io_masters_0_release_bits_header_src,
    output[1:0] io_masters_0_release_bits_header_dst,
    output[25:0] io_masters_0_release_bits_payload_addr,
    output[3:0] io_masters_0_release_bits_payload_client_xact_id,
    output[3:0] io_masters_0_release_bits_payload_master_xact_id,
    output[511:0] io_masters_0_release_bits_payload_data,
    output[2:0] io_masters_0_release_bits_payload_r_type
);

  wire T0;
  wire[3:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire[3:0] T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[511:0] T16;
  wire[1:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire[1:0] T23;
  wire[3:0] T24;
  wire[25:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire[1:0] T28;
  wire T29;
  wire T30;
  wire[2:0] T31;
  wire[511:0] T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire[25:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire T39;
  wire[2:0] T40;
  wire[511:0] T41;
  wire[3:0] T42;
  wire[3:0] T43;
  wire[25:0] T44;
  wire[1:0] T45;
  wire[1:0] T46;
  wire[1:0] T47;
  wire T48;
  wire T49;
  wire[3:0] T50;
  wire[2:0] T51;
  wire[5:0] T52;
  wire[2:0] T53;
  wire[511:0] T54;
  wire[3:0] T55;
  wire[25:0] T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire[3:0] T61;
  wire[2:0] T62;
  wire[5:0] T63;
  wire[2:0] T64;
  wire[511:0] T65;
  wire[3:0] T66;
  wire[25:0] T67;
  wire[1:0] T68;
  wire[1:0] T69;
  wire[1:0] T70;
  wire T71;
  wire[2:0] T72;
  wire[2:0] relNet_io_out_0_bits_payload_r_type;
  wire[511:0] T73;
  wire[511:0] relNet_io_out_0_bits_payload_data;
  wire[3:0] T74;
  wire[3:0] relNet_io_out_0_bits_payload_master_xact_id;
  wire[3:0] T75;
  wire[3:0] relNet_io_out_0_bits_payload_client_xact_id;
  wire[25:0] T76;
  wire[25:0] relNet_io_out_0_bits_payload_addr;
  wire[1:0] T77;
  wire[1:0] relNet_io_out_0_bits_header_dst;
  wire[1:0] T78;
  wire[1:0] T79;
  wire[1:0] relNet_io_out_0_bits_header_src;
  wire T80;
  wire relNet_io_out_0_valid;
  wire T81;
  wire prbNet_io_in_0_ready;
  wire[3:0] T82;
  wire[3:0] ackNet_io_out_0_bits_payload_master_xact_id;
  wire[1:0] T83;
  wire[1:0] ackNet_io_out_0_bits_header_dst;
  wire[1:0] T84;
  wire[1:0] T85;
  wire[1:0] ackNet_io_out_0_bits_header_src;
  wire T86;
  wire ackNet_io_out_0_valid;
  wire T87;
  wire gntNet_io_in_0_ready;
  wire[3:0] T88;
  wire[3:0] acqNet_io_out_0_bits_payload_atomic_opcode;
  wire[2:0] T89;
  wire[2:0] acqNet_io_out_0_bits_payload_subword_addr;
  wire[5:0] T90;
  wire[5:0] acqNet_io_out_0_bits_payload_write_mask;
  wire[2:0] T91;
  wire[2:0] acqNet_io_out_0_bits_payload_a_type;
  wire[511:0] T92;
  wire[511:0] acqNet_io_out_0_bits_payload_data;
  wire[3:0] T93;
  wire[3:0] acqNet_io_out_0_bits_payload_client_xact_id;
  wire[25:0] T94;
  wire[25:0] acqNet_io_out_0_bits_payload_addr;
  wire[1:0] T95;
  wire[1:0] acqNet_io_out_0_bits_header_dst;
  wire[1:0] T96;
  wire[1:0] T97;
  wire[1:0] acqNet_io_out_0_bits_header_src;
  wire T98;
  wire acqNet_io_out_0_valid;
  wire T99;
  wire relNet_io_in_1_ready;
  wire[1:0] T100;
  wire[1:0] prbNet_io_out_1_bits_payload_p_type;
  wire[3:0] T101;
  wire[3:0] prbNet_io_out_1_bits_payload_master_xact_id;
  wire[25:0] T102;
  wire[25:0] prbNet_io_out_1_bits_payload_addr;
  wire[1:0] T103;
  wire[1:0] T104;
  wire[1:0] prbNet_io_out_1_bits_header_dst;
  wire[1:0] T105;
  wire[1:0] prbNet_io_out_1_bits_header_src;
  wire T106;
  wire prbNet_io_out_1_valid;
  wire T107;
  wire ackNet_io_in_1_ready;
  wire[3:0] T108;
  wire[3:0] gntNet_io_out_1_bits_payload_g_type;
  wire[3:0] T109;
  wire[3:0] gntNet_io_out_1_bits_payload_master_xact_id;
  wire[3:0] T110;
  wire[3:0] gntNet_io_out_1_bits_payload_client_xact_id;
  wire[511:0] T111;
  wire[511:0] gntNet_io_out_1_bits_payload_data;
  wire[1:0] T112;
  wire[1:0] T113;
  wire[1:0] gntNet_io_out_1_bits_header_dst;
  wire[1:0] T114;
  wire[1:0] gntNet_io_out_1_bits_header_src;
  wire T115;
  wire gntNet_io_out_1_valid;
  wire T116;
  wire acqNet_io_in_1_ready;
  wire T117;
  wire relNet_io_in_2_ready;
  wire[1:0] T118;
  wire[1:0] prbNet_io_out_2_bits_payload_p_type;
  wire[3:0] T119;
  wire[3:0] prbNet_io_out_2_bits_payload_master_xact_id;
  wire[25:0] T120;
  wire[25:0] prbNet_io_out_2_bits_payload_addr;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] prbNet_io_out_2_bits_header_dst;
  wire[1:0] T123;
  wire[1:0] prbNet_io_out_2_bits_header_src;
  wire T124;
  wire prbNet_io_out_2_valid;
  wire T125;
  wire ackNet_io_in_2_ready;
  wire[3:0] T126;
  wire[3:0] gntNet_io_out_2_bits_payload_g_type;
  wire[3:0] T127;
  wire[3:0] gntNet_io_out_2_bits_payload_master_xact_id;
  wire[3:0] T128;
  wire[3:0] gntNet_io_out_2_bits_payload_client_xact_id;
  wire[511:0] T129;
  wire[511:0] gntNet_io_out_2_bits_payload_data;
  wire[1:0] T130;
  wire[1:0] T131;
  wire[1:0] gntNet_io_out_2_bits_header_dst;
  wire[1:0] T132;
  wire[1:0] gntNet_io_out_2_bits_header_src;
  wire T133;
  wire gntNet_io_out_2_valid;
  wire T134;
  wire acqNet_io_in_2_ready;


  assign T0 = io_masters_0_finish_ready;
  assign T1 = io_clients_0_finish_bits_payload_master_xact_id;
  assign T2 = io_clients_0_finish_bits_header_dst;
  assign T3 = T4;
  assign T4 = io_clients_0_finish_bits_header_src + 2'h1;
  assign T5 = io_clients_0_finish_valid;
  assign T6 = io_clients_1_finish_bits_payload_master_xact_id;
  assign T7 = io_clients_1_finish_bits_header_dst;
  assign T8 = T9;
  assign T9 = io_clients_1_finish_bits_header_src + 2'h1;
  assign T10 = io_clients_1_finish_valid;
  assign T11 = io_clients_0_grant_ready;
  assign T12 = io_clients_1_grant_ready;
  assign T13 = io_masters_0_grant_bits_payload_g_type;
  assign T14 = io_masters_0_grant_bits_payload_master_xact_id;
  assign T15 = io_masters_0_grant_bits_payload_client_xact_id;
  assign T16 = io_masters_0_grant_bits_payload_data;
  assign T17 = T18;
  assign T18 = io_masters_0_grant_bits_header_dst + 2'h1;
  assign T19 = io_masters_0_grant_bits_header_src;
  assign T20 = io_masters_0_grant_valid;
  assign T21 = io_clients_0_probe_ready;
  assign T22 = io_clients_1_probe_ready;
  assign T23 = io_masters_0_probe_bits_payload_p_type;
  assign T24 = io_masters_0_probe_bits_payload_master_xact_id;
  assign T25 = io_masters_0_probe_bits_payload_addr;
  assign T26 = T27;
  assign T27 = io_masters_0_probe_bits_header_dst + 2'h1;
  assign T28 = io_masters_0_probe_bits_header_src;
  assign T29 = io_masters_0_probe_valid;
  assign T30 = io_masters_0_release_ready;
  assign T31 = io_clients_0_release_bits_payload_r_type;
  assign T32 = io_clients_0_release_bits_payload_data;
  assign T33 = io_clients_0_release_bits_payload_master_xact_id;
  assign T34 = io_clients_0_release_bits_payload_client_xact_id;
  assign T35 = io_clients_0_release_bits_payload_addr;
  assign T36 = io_clients_0_release_bits_header_dst;
  assign T37 = T38;
  assign T38 = io_clients_0_release_bits_header_src + 2'h1;
  assign T39 = io_clients_0_release_valid;
  assign T40 = io_clients_1_release_bits_payload_r_type;
  assign T41 = io_clients_1_release_bits_payload_data;
  assign T42 = io_clients_1_release_bits_payload_master_xact_id;
  assign T43 = io_clients_1_release_bits_payload_client_xact_id;
  assign T44 = io_clients_1_release_bits_payload_addr;
  assign T45 = io_clients_1_release_bits_header_dst;
  assign T46 = T47;
  assign T47 = io_clients_1_release_bits_header_src + 2'h1;
  assign T48 = io_clients_1_release_valid;
  assign T49 = io_masters_0_acquire_ready;
  assign T50 = io_clients_0_acquire_bits_payload_atomic_opcode;
  assign T51 = io_clients_0_acquire_bits_payload_subword_addr;
  assign T52 = io_clients_0_acquire_bits_payload_write_mask;
  assign T53 = io_clients_0_acquire_bits_payload_a_type;
  assign T54 = io_clients_0_acquire_bits_payload_data;
  assign T55 = io_clients_0_acquire_bits_payload_client_xact_id;
  assign T56 = io_clients_0_acquire_bits_payload_addr;
  assign T57 = io_clients_0_acquire_bits_header_dst;
  assign T58 = T59;
  assign T59 = io_clients_0_acquire_bits_header_src + 2'h1;
  assign T60 = io_clients_0_acquire_valid;
  assign T61 = io_clients_1_acquire_bits_payload_atomic_opcode;
  assign T62 = io_clients_1_acquire_bits_payload_subword_addr;
  assign T63 = io_clients_1_acquire_bits_payload_write_mask;
  assign T64 = io_clients_1_acquire_bits_payload_a_type;
  assign T65 = io_clients_1_acquire_bits_payload_data;
  assign T66 = io_clients_1_acquire_bits_payload_client_xact_id;
  assign T67 = io_clients_1_acquire_bits_payload_addr;
  assign T68 = io_clients_1_acquire_bits_header_dst;
  assign T69 = T70;
  assign T70 = io_clients_1_acquire_bits_header_src + 2'h1;
  assign T71 = io_clients_1_acquire_valid;
  assign io_masters_0_release_bits_payload_r_type = T72;
  assign T72 = relNet_io_out_0_bits_payload_r_type;
  assign io_masters_0_release_bits_payload_data = T73;
  assign T73 = relNet_io_out_0_bits_payload_data;
  assign io_masters_0_release_bits_payload_master_xact_id = T74;
  assign T74 = relNet_io_out_0_bits_payload_master_xact_id;
  assign io_masters_0_release_bits_payload_client_xact_id = T75;
  assign T75 = relNet_io_out_0_bits_payload_client_xact_id;
  assign io_masters_0_release_bits_payload_addr = T76;
  assign T76 = relNet_io_out_0_bits_payload_addr;
  assign io_masters_0_release_bits_header_dst = T77;
  assign T77 = relNet_io_out_0_bits_header_dst;
  assign io_masters_0_release_bits_header_src = T78;
  assign T78 = T79;
  assign T79 = relNet_io_out_0_bits_header_src - 2'h1;
  assign io_masters_0_release_valid = T80;
  assign T80 = relNet_io_out_0_valid;
  assign io_masters_0_probe_ready = T81;
  assign T81 = prbNet_io_in_0_ready;
  assign io_masters_0_finish_bits_payload_master_xact_id = T82;
  assign T82 = ackNet_io_out_0_bits_payload_master_xact_id;
  assign io_masters_0_finish_bits_header_dst = T83;
  assign T83 = ackNet_io_out_0_bits_header_dst;
  assign io_masters_0_finish_bits_header_src = T84;
  assign T84 = T85;
  assign T85 = ackNet_io_out_0_bits_header_src - 2'h1;
  assign io_masters_0_finish_valid = T86;
  assign T86 = ackNet_io_out_0_valid;
  assign io_masters_0_grant_ready = T87;
  assign T87 = gntNet_io_in_0_ready;
  assign io_masters_0_acquire_bits_payload_atomic_opcode = T88;
  assign T88 = acqNet_io_out_0_bits_payload_atomic_opcode;
  assign io_masters_0_acquire_bits_payload_subword_addr = T89;
  assign T89 = acqNet_io_out_0_bits_payload_subword_addr;
  assign io_masters_0_acquire_bits_payload_write_mask = T90;
  assign T90 = acqNet_io_out_0_bits_payload_write_mask;
  assign io_masters_0_acquire_bits_payload_a_type = T91;
  assign T91 = acqNet_io_out_0_bits_payload_a_type;
  assign io_masters_0_acquire_bits_payload_data = T92;
  assign T92 = acqNet_io_out_0_bits_payload_data;
  assign io_masters_0_acquire_bits_payload_client_xact_id = T93;
  assign T93 = acqNet_io_out_0_bits_payload_client_xact_id;
  assign io_masters_0_acquire_bits_payload_addr = T94;
  assign T94 = acqNet_io_out_0_bits_payload_addr;
  assign io_masters_0_acquire_bits_header_dst = T95;
  assign T95 = acqNet_io_out_0_bits_header_dst;
  assign io_masters_0_acquire_bits_header_src = T96;
  assign T96 = T97;
  assign T97 = acqNet_io_out_0_bits_header_src - 2'h1;
  assign io_masters_0_acquire_valid = T98;
  assign T98 = acqNet_io_out_0_valid;
  assign io_clients_0_release_ready = T99;
  assign T99 = relNet_io_in_1_ready;
  assign io_clients_0_probe_bits_payload_p_type = T100;
  assign T100 = prbNet_io_out_1_bits_payload_p_type;
  assign io_clients_0_probe_bits_payload_master_xact_id = T101;
  assign T101 = prbNet_io_out_1_bits_payload_master_xact_id;
  assign io_clients_0_probe_bits_payload_addr = T102;
  assign T102 = prbNet_io_out_1_bits_payload_addr;
  assign io_clients_0_probe_bits_header_dst = T103;
  assign T103 = T104;
  assign T104 = prbNet_io_out_1_bits_header_dst - 2'h1;
  assign io_clients_0_probe_bits_header_src = T105;
  assign T105 = prbNet_io_out_1_bits_header_src;
  assign io_clients_0_probe_valid = T106;
  assign T106 = prbNet_io_out_1_valid;
  assign io_clients_0_finish_ready = T107;
  assign T107 = ackNet_io_in_1_ready;
  assign io_clients_0_grant_bits_payload_g_type = T108;
  assign T108 = gntNet_io_out_1_bits_payload_g_type;
  assign io_clients_0_grant_bits_payload_master_xact_id = T109;
  assign T109 = gntNet_io_out_1_bits_payload_master_xact_id;
  assign io_clients_0_grant_bits_payload_client_xact_id = T110;
  assign T110 = gntNet_io_out_1_bits_payload_client_xact_id;
  assign io_clients_0_grant_bits_payload_data = T111;
  assign T111 = gntNet_io_out_1_bits_payload_data;
  assign io_clients_0_grant_bits_header_dst = T112;
  assign T112 = T113;
  assign T113 = gntNet_io_out_1_bits_header_dst - 2'h1;
  assign io_clients_0_grant_bits_header_src = T114;
  assign T114 = gntNet_io_out_1_bits_header_src;
  assign io_clients_0_grant_valid = T115;
  assign T115 = gntNet_io_out_1_valid;
  assign io_clients_0_acquire_ready = T116;
  assign T116 = acqNet_io_in_1_ready;
  assign io_clients_1_release_ready = T117;
  assign T117 = relNet_io_in_2_ready;
  assign io_clients_1_probe_bits_payload_p_type = T118;
  assign T118 = prbNet_io_out_2_bits_payload_p_type;
  assign io_clients_1_probe_bits_payload_master_xact_id = T119;
  assign T119 = prbNet_io_out_2_bits_payload_master_xact_id;
  assign io_clients_1_probe_bits_payload_addr = T120;
  assign T120 = prbNet_io_out_2_bits_payload_addr;
  assign io_clients_1_probe_bits_header_dst = T121;
  assign T121 = T122;
  assign T122 = prbNet_io_out_2_bits_header_dst - 2'h1;
  assign io_clients_1_probe_bits_header_src = T123;
  assign T123 = prbNet_io_out_2_bits_header_src;
  assign io_clients_1_probe_valid = T124;
  assign T124 = prbNet_io_out_2_valid;
  assign io_clients_1_finish_ready = T125;
  assign T125 = ackNet_io_in_2_ready;
  assign io_clients_1_grant_bits_payload_g_type = T126;
  assign T126 = gntNet_io_out_2_bits_payload_g_type;
  assign io_clients_1_grant_bits_payload_master_xact_id = T127;
  assign T127 = gntNet_io_out_2_bits_payload_master_xact_id;
  assign io_clients_1_grant_bits_payload_client_xact_id = T128;
  assign T128 = gntNet_io_out_2_bits_payload_client_xact_id;
  assign io_clients_1_grant_bits_payload_data = T129;
  assign T129 = gntNet_io_out_2_bits_payload_data;
  assign io_clients_1_grant_bits_header_dst = T130;
  assign T130 = T131;
  assign T131 = gntNet_io_out_2_bits_header_dst - 2'h1;
  assign io_clients_1_grant_bits_header_src = T132;
  assign T132 = gntNet_io_out_2_bits_header_src;
  assign io_clients_1_grant_valid = T133;
  assign T133 = gntNet_io_out_2_valid;
  assign io_clients_1_acquire_ready = T134;
  assign T134 = acqNet_io_in_2_ready;
  BasicCrossbar_0 acqNet(.clk(clk), .reset(reset),
       .io_in_2_ready( acqNet_io_in_2_ready ),
       .io_in_2_valid( T71 ),
       .io_in_2_bits_header_src( T69 ),
       .io_in_2_bits_header_dst( T68 ),
       .io_in_2_bits_payload_addr( T67 ),
       .io_in_2_bits_payload_client_xact_id( T66 ),
       .io_in_2_bits_payload_data( T65 ),
       .io_in_2_bits_payload_a_type( T64 ),
       .io_in_2_bits_payload_write_mask( T63 ),
       .io_in_2_bits_payload_subword_addr( T62 ),
       .io_in_2_bits_payload_atomic_opcode( T61 ),
       .io_in_1_ready( acqNet_io_in_1_ready ),
       .io_in_1_valid( T60 ),
       .io_in_1_bits_header_src( T58 ),
       .io_in_1_bits_header_dst( T57 ),
       .io_in_1_bits_payload_addr( T56 ),
       .io_in_1_bits_payload_client_xact_id( T55 ),
       .io_in_1_bits_payload_data( T54 ),
       .io_in_1_bits_payload_a_type( T53 ),
       .io_in_1_bits_payload_write_mask( T52 ),
       .io_in_1_bits_payload_subword_addr( T51 ),
       .io_in_1_bits_payload_atomic_opcode( T50 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_client_xact_id(  )
       //.io_in_0_bits_payload_data(  )
       //.io_in_0_bits_payload_a_type(  )
       //.io_in_0_bits_payload_write_mask(  )
       //.io_in_0_bits_payload_subword_addr(  )
       //.io_in_0_bits_payload_atomic_opcode(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_addr(  )
       //.io_out_2_bits_payload_client_xact_id(  )
       //.io_out_2_bits_payload_data(  )
       //.io_out_2_bits_payload_a_type(  )
       //.io_out_2_bits_payload_write_mask(  )
       //.io_out_2_bits_payload_subword_addr(  )
       //.io_out_2_bits_payload_atomic_opcode(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_addr(  )
       //.io_out_1_bits_payload_client_xact_id(  )
       //.io_out_1_bits_payload_data(  )
       //.io_out_1_bits_payload_a_type(  )
       //.io_out_1_bits_payload_write_mask(  )
       //.io_out_1_bits_payload_subword_addr(  )
       //.io_out_1_bits_payload_atomic_opcode(  )
       .io_out_0_ready( T49 ),
       .io_out_0_valid( acqNet_io_out_0_valid ),
       .io_out_0_bits_header_src( acqNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( acqNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_addr( acqNet_io_out_0_bits_payload_addr ),
       .io_out_0_bits_payload_client_xact_id( acqNet_io_out_0_bits_payload_client_xact_id ),
       .io_out_0_bits_payload_data( acqNet_io_out_0_bits_payload_data ),
       .io_out_0_bits_payload_a_type( acqNet_io_out_0_bits_payload_a_type ),
       .io_out_0_bits_payload_write_mask( acqNet_io_out_0_bits_payload_write_mask ),
       .io_out_0_bits_payload_subword_addr( acqNet_io_out_0_bits_payload_subword_addr ),
       .io_out_0_bits_payload_atomic_opcode( acqNet_io_out_0_bits_payload_atomic_opcode )
  );
  `ifndef SYNTHESIS
    assign acqNet.io_in_0_bits_header_src = {1{$random}};
    assign acqNet.io_in_0_bits_header_dst = {1{$random}};
    assign acqNet.io_in_0_bits_payload_addr = {1{$random}};
    assign acqNet.io_in_0_bits_payload_client_xact_id = {1{$random}};
    assign acqNet.io_in_0_bits_payload_data = {16{$random}};
    assign acqNet.io_in_0_bits_payload_a_type = {1{$random}};
    assign acqNet.io_in_0_bits_payload_write_mask = {1{$random}};
    assign acqNet.io_in_0_bits_payload_subword_addr = {1{$random}};
    assign acqNet.io_in_0_bits_payload_atomic_opcode = {1{$random}};
  `endif
  BasicCrossbar_1 relNet(.clk(clk), .reset(reset),
       .io_in_2_ready( relNet_io_in_2_ready ),
       .io_in_2_valid( T48 ),
       .io_in_2_bits_header_src( T46 ),
       .io_in_2_bits_header_dst( T45 ),
       .io_in_2_bits_payload_addr( T44 ),
       .io_in_2_bits_payload_client_xact_id( T43 ),
       .io_in_2_bits_payload_master_xact_id( T42 ),
       .io_in_2_bits_payload_data( T41 ),
       .io_in_2_bits_payload_r_type( T40 ),
       .io_in_1_ready( relNet_io_in_1_ready ),
       .io_in_1_valid( T39 ),
       .io_in_1_bits_header_src( T37 ),
       .io_in_1_bits_header_dst( T36 ),
       .io_in_1_bits_payload_addr( T35 ),
       .io_in_1_bits_payload_client_xact_id( T34 ),
       .io_in_1_bits_payload_master_xact_id( T33 ),
       .io_in_1_bits_payload_data( T32 ),
       .io_in_1_bits_payload_r_type( T31 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_client_xact_id(  )
       //.io_in_0_bits_payload_master_xact_id(  )
       //.io_in_0_bits_payload_data(  )
       //.io_in_0_bits_payload_r_type(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_addr(  )
       //.io_out_2_bits_payload_client_xact_id(  )
       //.io_out_2_bits_payload_master_xact_id(  )
       //.io_out_2_bits_payload_data(  )
       //.io_out_2_bits_payload_r_type(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_addr(  )
       //.io_out_1_bits_payload_client_xact_id(  )
       //.io_out_1_bits_payload_master_xact_id(  )
       //.io_out_1_bits_payload_data(  )
       //.io_out_1_bits_payload_r_type(  )
       .io_out_0_ready( T30 ),
       .io_out_0_valid( relNet_io_out_0_valid ),
       .io_out_0_bits_header_src( relNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( relNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_addr( relNet_io_out_0_bits_payload_addr ),
       .io_out_0_bits_payload_client_xact_id( relNet_io_out_0_bits_payload_client_xact_id ),
       .io_out_0_bits_payload_master_xact_id( relNet_io_out_0_bits_payload_master_xact_id ),
       .io_out_0_bits_payload_data( relNet_io_out_0_bits_payload_data ),
       .io_out_0_bits_payload_r_type( relNet_io_out_0_bits_payload_r_type )
  );
  `ifndef SYNTHESIS
    assign relNet.io_in_0_bits_header_src = {1{$random}};
    assign relNet.io_in_0_bits_header_dst = {1{$random}};
    assign relNet.io_in_0_bits_payload_addr = {1{$random}};
    assign relNet.io_in_0_bits_payload_client_xact_id = {1{$random}};
    assign relNet.io_in_0_bits_payload_master_xact_id = {1{$random}};
    assign relNet.io_in_0_bits_payload_data = {16{$random}};
    assign relNet.io_in_0_bits_payload_r_type = {1{$random}};
  `endif
  BasicCrossbar_2 prbNet(.clk(clk), .reset(reset),
       //.io_in_2_ready(  )
       .io_in_2_valid( 1'h0 ),
       //.io_in_2_bits_header_src(  )
       //.io_in_2_bits_header_dst(  )
       //.io_in_2_bits_payload_addr(  )
       //.io_in_2_bits_payload_master_xact_id(  )
       //.io_in_2_bits_payload_p_type(  )
       //.io_in_1_ready(  )
       .io_in_1_valid( 1'h0 ),
       //.io_in_1_bits_header_src(  )
       //.io_in_1_bits_header_dst(  )
       //.io_in_1_bits_payload_addr(  )
       //.io_in_1_bits_payload_master_xact_id(  )
       //.io_in_1_bits_payload_p_type(  )
       .io_in_0_ready( prbNet_io_in_0_ready ),
       .io_in_0_valid( T29 ),
       .io_in_0_bits_header_src( T28 ),
       .io_in_0_bits_header_dst( T26 ),
       .io_in_0_bits_payload_addr( T25 ),
       .io_in_0_bits_payload_master_xact_id( T24 ),
       .io_in_0_bits_payload_p_type( T23 ),
       .io_out_2_ready( T22 ),
       .io_out_2_valid( prbNet_io_out_2_valid ),
       .io_out_2_bits_header_src( prbNet_io_out_2_bits_header_src ),
       .io_out_2_bits_header_dst( prbNet_io_out_2_bits_header_dst ),
       .io_out_2_bits_payload_addr( prbNet_io_out_2_bits_payload_addr ),
       .io_out_2_bits_payload_master_xact_id( prbNet_io_out_2_bits_payload_master_xact_id ),
       .io_out_2_bits_payload_p_type( prbNet_io_out_2_bits_payload_p_type ),
       .io_out_1_ready( T21 ),
       .io_out_1_valid( prbNet_io_out_1_valid ),
       .io_out_1_bits_header_src( prbNet_io_out_1_bits_header_src ),
       .io_out_1_bits_header_dst( prbNet_io_out_1_bits_header_dst ),
       .io_out_1_bits_payload_addr( prbNet_io_out_1_bits_payload_addr ),
       .io_out_1_bits_payload_master_xact_id( prbNet_io_out_1_bits_payload_master_xact_id ),
       .io_out_1_bits_payload_p_type( prbNet_io_out_1_bits_payload_p_type ),
       .io_out_0_ready( 1'h0 )
       //.io_out_0_valid(  )
       //.io_out_0_bits_header_src(  )
       //.io_out_0_bits_header_dst(  )
       //.io_out_0_bits_payload_addr(  )
       //.io_out_0_bits_payload_master_xact_id(  )
       //.io_out_0_bits_payload_p_type(  )
  );
  `ifndef SYNTHESIS
    assign prbNet.io_in_2_bits_header_src = {1{$random}};
    assign prbNet.io_in_2_bits_header_dst = {1{$random}};
    assign prbNet.io_in_2_bits_payload_addr = {1{$random}};
    assign prbNet.io_in_2_bits_payload_master_xact_id = {1{$random}};
    assign prbNet.io_in_2_bits_payload_p_type = {1{$random}};
    assign prbNet.io_in_1_bits_header_src = {1{$random}};
    assign prbNet.io_in_1_bits_header_dst = {1{$random}};
    assign prbNet.io_in_1_bits_payload_addr = {1{$random}};
    assign prbNet.io_in_1_bits_payload_master_xact_id = {1{$random}};
    assign prbNet.io_in_1_bits_payload_p_type = {1{$random}};
  `endif
  BasicCrossbar_3 gntNet(.clk(clk), .reset(reset),
       //.io_in_2_ready(  )
       .io_in_2_valid( 1'h0 ),
       //.io_in_2_bits_header_src(  )
       //.io_in_2_bits_header_dst(  )
       //.io_in_2_bits_payload_data(  )
       //.io_in_2_bits_payload_client_xact_id(  )
       //.io_in_2_bits_payload_master_xact_id(  )
       //.io_in_2_bits_payload_g_type(  )
       //.io_in_1_ready(  )
       .io_in_1_valid( 1'h0 ),
       //.io_in_1_bits_header_src(  )
       //.io_in_1_bits_header_dst(  )
       //.io_in_1_bits_payload_data(  )
       //.io_in_1_bits_payload_client_xact_id(  )
       //.io_in_1_bits_payload_master_xact_id(  )
       //.io_in_1_bits_payload_g_type(  )
       .io_in_0_ready( gntNet_io_in_0_ready ),
       .io_in_0_valid( T20 ),
       .io_in_0_bits_header_src( T19 ),
       .io_in_0_bits_header_dst( T17 ),
       .io_in_0_bits_payload_data( T16 ),
       .io_in_0_bits_payload_client_xact_id( T15 ),
       .io_in_0_bits_payload_master_xact_id( T14 ),
       .io_in_0_bits_payload_g_type( T13 ),
       .io_out_2_ready( T12 ),
       .io_out_2_valid( gntNet_io_out_2_valid ),
       .io_out_2_bits_header_src( gntNet_io_out_2_bits_header_src ),
       .io_out_2_bits_header_dst( gntNet_io_out_2_bits_header_dst ),
       .io_out_2_bits_payload_data( gntNet_io_out_2_bits_payload_data ),
       .io_out_2_bits_payload_client_xact_id( gntNet_io_out_2_bits_payload_client_xact_id ),
       .io_out_2_bits_payload_master_xact_id( gntNet_io_out_2_bits_payload_master_xact_id ),
       .io_out_2_bits_payload_g_type( gntNet_io_out_2_bits_payload_g_type ),
       .io_out_1_ready( T11 ),
       .io_out_1_valid( gntNet_io_out_1_valid ),
       .io_out_1_bits_header_src( gntNet_io_out_1_bits_header_src ),
       .io_out_1_bits_header_dst( gntNet_io_out_1_bits_header_dst ),
       .io_out_1_bits_payload_data( gntNet_io_out_1_bits_payload_data ),
       .io_out_1_bits_payload_client_xact_id( gntNet_io_out_1_bits_payload_client_xact_id ),
       .io_out_1_bits_payload_master_xact_id( gntNet_io_out_1_bits_payload_master_xact_id ),
       .io_out_1_bits_payload_g_type( gntNet_io_out_1_bits_payload_g_type ),
       .io_out_0_ready( 1'h0 )
       //.io_out_0_valid(  )
       //.io_out_0_bits_header_src(  )
       //.io_out_0_bits_header_dst(  )
       //.io_out_0_bits_payload_data(  )
       //.io_out_0_bits_payload_client_xact_id(  )
       //.io_out_0_bits_payload_master_xact_id(  )
       //.io_out_0_bits_payload_g_type(  )
  );
  `ifndef SYNTHESIS
    assign gntNet.io_in_2_bits_header_src = {1{$random}};
    assign gntNet.io_in_2_bits_header_dst = {1{$random}};
    assign gntNet.io_in_2_bits_payload_data = {16{$random}};
    assign gntNet.io_in_2_bits_payload_client_xact_id = {1{$random}};
    assign gntNet.io_in_2_bits_payload_master_xact_id = {1{$random}};
    assign gntNet.io_in_2_bits_payload_g_type = {1{$random}};
    assign gntNet.io_in_1_bits_header_src = {1{$random}};
    assign gntNet.io_in_1_bits_header_dst = {1{$random}};
    assign gntNet.io_in_1_bits_payload_data = {16{$random}};
    assign gntNet.io_in_1_bits_payload_client_xact_id = {1{$random}};
    assign gntNet.io_in_1_bits_payload_master_xact_id = {1{$random}};
    assign gntNet.io_in_1_bits_payload_g_type = {1{$random}};
  `endif
  BasicCrossbar_4 ackNet(.clk(clk), .reset(reset),
       .io_in_2_ready( ackNet_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( T8 ),
       .io_in_2_bits_header_dst( T7 ),
       .io_in_2_bits_payload_master_xact_id( T6 ),
       .io_in_1_ready( ackNet_io_in_1_ready ),
       .io_in_1_valid( T5 ),
       .io_in_1_bits_header_src( T3 ),
       .io_in_1_bits_header_dst( T2 ),
       .io_in_1_bits_payload_master_xact_id( T1 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_master_xact_id(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_master_xact_id(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_master_xact_id(  )
       .io_out_0_ready( T0 ),
       .io_out_0_valid( ackNet_io_out_0_valid ),
       .io_out_0_bits_header_src( ackNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( ackNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_master_xact_id( ackNet_io_out_0_bits_payload_master_xact_id )
  );
  `ifndef SYNTHESIS
    assign ackNet.io_in_0_bits_header_src = {1{$random}};
    assign ackNet.io_in_0_bits_header_dst = {1{$random}};
    assign ackNet.io_in_0_bits_payload_master_xact_id = {1{$random}};
  `endif
endmodule

module Queue_3(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [4:0] io_enq_bits_tag,
    input  io_enq_bits_rw,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[4:0] io_deq_bits_tag,
    output io_deq_bits_rw,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  deq_ptr;
  wire T1;
  wire T2;
  wire T3;
  wire do_deq;
  wire T4;
  wire do_flow;
  wire T5;
  reg  enq_ptr;
  wire T6;
  wire T7;
  wire T8;
  wire do_enq;
  wire T9;
  wire T10;
  wire T11;
  wire ptr_match;
  reg  maybe_full;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[31:0] T16;
  wire[5:0] T17;
  wire T18;
  wire[31:0] T19;
  reg [31:0] ram [1:0];
  wire[31:0] T20;
  wire[31:0] T21;
  wire[31:0] T22;
  wire[5:0] T23;
  wire[4:0] T24;
  wire[25:0] T25;
  wire[4:0] T26;
  wire[25:0] T27;
  wire T28;
  wire empty;
  wire T29;
  wire T30;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    deq_ptr = {1{$random}};
    enq_ptr = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T11, ptr_diff};
  assign ptr_diff = enq_ptr - deq_ptr;
  assign T1 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : deq_ptr;
  assign T3 = deq_ptr + 1'h1;
  assign do_deq = T5 & T4;
  assign T4 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T5 = io_deq_ready & io_deq_valid;
  assign T6 = reset ? 1'h0 : T7;
  assign T7 = do_enq ? T8 : enq_ptr;
  assign T8 = enq_ptr + 1'h1;
  assign do_enq = T10 & T9;
  assign T9 = do_flow ^ 1'h1;
  assign T10 = io_enq_ready & io_enq_valid;
  assign T11 = maybe_full & ptr_match;
  assign ptr_match = enq_ptr == deq_ptr;
  assign T12 = reset ? 1'h0 : T13;
  assign T13 = T14 ? do_enq : maybe_full;
  assign T14 = do_enq != do_deq;
  assign io_deq_bits_rw = T15;
  assign T15 = T16[1'h0:1'h0];
  assign T16 = {T25, T17};
  assign T17 = {T24, T18};
  assign T18 = T19[1'h0:1'h0];
  assign T19 = ram[deq_ptr];
  always @(posedge clk)
    if (do_enq)
      ram[enq_ptr] <= T21;
  assign T21 = T22;
  assign T22 = {io_enq_bits_addr, T23};
  assign T23 = {io_enq_bits_tag, io_enq_bits_rw};
  assign T24 = T19[3'h5:1'h1];
  assign T25 = T19[5'h1f:3'h6];
  assign io_deq_bits_tag = T26;
  assign T26 = T16[3'h5:1'h1];
  assign io_deq_bits_addr = T27;
  assign T27 = T16[5'h1f:3'h6];
  assign io_deq_valid = T28;
  assign T28 = empty ^ 1'h1;
  assign empty = ptr_match & T29;
  assign T29 = maybe_full ^ 1'h1;
  assign io_enq_ready = T30;
  assign T30 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      deq_ptr <= 1'h0;
    end else if(do_deq) begin
      deq_ptr <= T3;
    end
    if(reset) begin
      enq_ptr <= 1'h0;
    end else if(do_enq) begin
      enq_ptr <= T8;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T14) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_4(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  deq_ptr;
  wire T1;
  wire T2;
  wire T3;
  wire do_deq;
  wire T4;
  wire do_flow;
  wire T5;
  reg  enq_ptr;
  wire T6;
  wire T7;
  wire T8;
  wire do_enq;
  wire T9;
  wire T10;
  wire T11;
  wire ptr_match;
  reg  maybe_full;
  wire T12;
  wire T13;
  wire T14;
  wire[127:0] T15;
  wire[127:0] T16;
  reg [127:0] ram [1:0];
  wire[127:0] T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    deq_ptr = {1{$random}};
    enq_ptr = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {4{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T11, ptr_diff};
  assign ptr_diff = enq_ptr - deq_ptr;
  assign T1 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : deq_ptr;
  assign T3 = deq_ptr + 1'h1;
  assign do_deq = T5 & T4;
  assign T4 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T5 = io_deq_ready & io_deq_valid;
  assign T6 = reset ? 1'h0 : T7;
  assign T7 = do_enq ? T8 : enq_ptr;
  assign T8 = enq_ptr + 1'h1;
  assign do_enq = T10 & T9;
  assign T9 = do_flow ^ 1'h1;
  assign T10 = io_enq_ready & io_enq_valid;
  assign T11 = maybe_full & ptr_match;
  assign ptr_match = enq_ptr == deq_ptr;
  assign T12 = reset ? 1'h0 : T13;
  assign T13 = T14 ? do_enq : maybe_full;
  assign T14 = do_enq != do_deq;
  assign io_deq_bits_data = T15;
  assign T15 = T16[7'h7f:1'h0];
  assign T16 = ram[deq_ptr];
  always @(posedge clk)
    if (do_enq)
      ram[enq_ptr] <= io_enq_bits_data;
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      deq_ptr <= 1'h0;
    end else if(do_deq) begin
      deq_ptr <= T3;
    end
    if(reset) begin
      enq_ptr <= 1'h0;
    end else if(do_enq) begin
      enq_ptr <= T8;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T14) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module MemIOUncachedTileLinkIOConverter(input clk, input reset,
    output io_uncached_acquire_ready,
    input  io_uncached_acquire_valid,
    input [1:0] io_uncached_acquire_bits_header_src,
    input [1:0] io_uncached_acquire_bits_header_dst,
    input [25:0] io_uncached_acquire_bits_payload_addr,
    input [3:0] io_uncached_acquire_bits_payload_client_xact_id,
    input [511:0] io_uncached_acquire_bits_payload_data,
    input [2:0] io_uncached_acquire_bits_payload_a_type,
    input [5:0] io_uncached_acquire_bits_payload_write_mask,
    input [2:0] io_uncached_acquire_bits_payload_subword_addr,
    input [3:0] io_uncached_acquire_bits_payload_atomic_opcode,
    input  io_uncached_grant_ready,
    output io_uncached_grant_valid,
    //output[1:0] io_uncached_grant_bits_header_src
    //output[1:0] io_uncached_grant_bits_header_dst
    output[511:0] io_uncached_grant_bits_payload_data,
    output[3:0] io_uncached_grant_bits_payload_client_xact_id,
    output[3:0] io_uncached_grant_bits_payload_master_xact_id,
    output[3:0] io_uncached_grant_bits_payload_g_type,
    //output io_uncached_finish_ready
    input  io_uncached_finish_valid,
    input [1:0] io_uncached_finish_bits_header_src,
    input [1:0] io_uncached_finish_bits_header_dst,
    input [3:0] io_uncached_finish_bits_payload_master_xact_id,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    output io_mem_resp_ready,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
);

  wire[127:0] T0;
  reg [511:0] buf_out;
  wire[511:0] T1;
  wire[511:0] T2;
  wire T3;
  wire T4;
  reg  active_out;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  reg [2:0] cnt_out;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire T15;
  wire T16;
  wire mem_data_q_io_enq_ready;
  wire T17;
  reg  has_data;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  reg  cmd_sent_out;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire mem_cmd_q_io_enq_ready;
  wire[511:0] T30;
  wire[383:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire[4:0] T35;
  reg [3:0] tag_out;
  wire[3:0] T36;
  reg [25:0] addr_out;
  wire[25:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  reg [2:0] cnt_in;
  wire[2:0] T42;
  wire[2:0] T43;
  wire T44;
  wire T45;
  reg  active_in;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[2:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire[127:0] mem_data_q_io_deq_bits_data;
  wire mem_data_q_io_deq_valid;
  wire mem_cmd_q_io_deq_bits_rw;
  wire[4:0] mem_cmd_q_io_deq_bits_tag;
  wire[25:0] mem_cmd_q_io_deq_bits_addr;
  wire mem_cmd_q_io_deq_valid;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] T57;
  wire[3:0] T58;
  reg [4:0] tag_in;
  wire[4:0] T59;
  wire[511:0] T60;
  reg [511:0] buf_in;
  wire[511:0] T61;
  wire[511:0] T62;
  wire[511:0] T63;
  wire[511:0] T64;
  wire[383:0] T65;
  wire T66;
  wire T67;
  wire T68;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    buf_out = {16{$random}};
    active_out = {1{$random}};
    cnt_out = {1{$random}};
    has_data = {1{$random}};
    cmd_sent_out = {1{$random}};
    tag_out = {1{$random}};
    addr_out = {1{$random}};
    cnt_in = {1{$random}};
    active_in = {1{$random}};
    tag_in = {1{$random}};
    buf_in = {16{$random}};
  end
`endif

  assign T0 = buf_out[7'h7f:1'h0];
  assign T1 = T15 ? T30 : T2;
  assign T2 = T3 ? io_uncached_acquire_bits_payload_data : buf_out;
  assign T3 = T4 & io_uncached_acquire_valid;
  assign T4 = active_out ^ 1'h1;
  assign T5 = reset ? 1'h0 : T6;
  assign T6 = T8 ? 1'h0 : T7;
  assign T7 = T3 ? 1'h1 : active_out;
  assign T8 = active_out & T9;
  assign T9 = cmd_sent_out & T10;
  assign T10 = T17 | T11;
  assign T11 = cnt_out == 3'h4;
  assign T12 = T15 ? T14 : T13;
  assign T13 = T3 ? 3'h0 : cnt_out;
  assign T14 = cnt_out + 3'h1;
  assign T15 = active_out & T16;
  assign T16 = mem_data_q_io_enq_ready & T32;
  assign T17 = has_data ^ 1'h1;
  assign T18 = reset ? 1'h0 : T19;
  assign T19 = T3 ? T20 : has_data;
  assign T20 = T22 | T21;
  assign T21 = 3'h6 == io_uncached_acquire_bits_payload_a_type;
  assign T22 = T24 | T23;
  assign T23 = 3'h5 == io_uncached_acquire_bits_payload_a_type;
  assign T24 = 3'h3 == io_uncached_acquire_bits_payload_a_type;
  assign T25 = reset ? 1'h0 : T26;
  assign T26 = T28 ? 1'h1 : T27;
  assign T27 = T3 ? 1'h0 : cmd_sent_out;
  assign T28 = active_out & T29;
  assign T29 = mem_cmd_q_io_enq_ready & T38;
  assign T30 = {128'h0, T31};
  assign T31 = buf_out >> 8'h80;
  assign T32 = T34 & T33;
  assign T33 = cnt_out < 3'h4;
  assign T34 = active_out & has_data;
  assign T35 = {1'h0, tag_out};
  assign T36 = T3 ? io_uncached_acquire_bits_payload_client_xact_id : tag_out;
  assign T37 = T3 ? io_uncached_acquire_bits_payload_addr : addr_out;
  assign T38 = active_out & T39;
  assign T39 = cmd_sent_out ^ 1'h1;
  assign io_mem_resp_ready = T40;
  assign T40 = T54 | T41;
  assign T41 = cnt_in < 3'h4;
  assign T42 = T52 ? T51 : T43;
  assign T43 = T44 ? 3'h1 : cnt_in;
  assign T44 = T45 & io_mem_resp_valid;
  assign T45 = active_in ^ 1'h1;
  assign T46 = reset ? 1'h0 : T47;
  assign T47 = T49 ? 1'h0 : T48;
  assign T48 = T44 ? 1'h1 : active_in;
  assign T49 = active_in & T50;
  assign T50 = io_uncached_grant_ready & io_uncached_grant_valid;
  assign T51 = cnt_in + 3'h1;
  assign T52 = active_in & T53;
  assign T53 = io_mem_resp_ready & io_mem_resp_valid;
  assign T54 = active_in ^ 1'h1;
  assign io_mem_req_data_bits_data = mem_data_q_io_deq_bits_data;
  assign io_mem_req_data_valid = mem_data_q_io_deq_valid;
  assign io_mem_req_cmd_bits_rw = mem_cmd_q_io_deq_bits_rw;
  assign io_mem_req_cmd_bits_tag = mem_cmd_q_io_deq_bits_tag;
  assign io_mem_req_cmd_bits_addr = mem_cmd_q_io_deq_bits_addr;
  assign io_mem_req_cmd_valid = mem_cmd_q_io_deq_valid;
  assign io_uncached_grant_bits_payload_g_type = T55;
  assign T55 = 4'h0;
  assign io_uncached_grant_bits_payload_master_xact_id = T56;
  assign T56 = 4'h0;
  assign io_uncached_grant_bits_payload_client_xact_id = T57;
  assign T57 = T58;
  assign T58 = tag_in[2'h3:1'h0];
  assign T59 = T44 ? io_mem_resp_bits_tag : tag_in;
  assign io_uncached_grant_bits_payload_data = T60;
  assign T60 = buf_in;
  assign T61 = T52 ? T64 : T62;
  assign T62 = T44 ? T63 : buf_in;
  assign T63 = io_mem_resp_bits_data << 9'h180;
  assign T64 = {io_mem_resp_bits_data, T65};
  assign T65 = buf_in[9'h1ff:8'h80];
  assign io_uncached_grant_valid = T66;
  assign T66 = active_in & T67;
  assign T67 = cnt_in == 3'h4;
  assign io_uncached_acquire_ready = T68;
  assign T68 = active_out ^ 1'h1;
  Queue_3 mem_cmd_q(.clk(clk), .reset(reset),
       .io_enq_ready( mem_cmd_q_io_enq_ready ),
       .io_enq_valid( T38 ),
       .io_enq_bits_addr( addr_out ),
       .io_enq_bits_tag( T35 ),
       .io_enq_bits_rw( has_data ),
       .io_deq_ready( io_mem_req_cmd_ready ),
       .io_deq_valid( mem_cmd_q_io_deq_valid ),
       .io_deq_bits_addr( mem_cmd_q_io_deq_bits_addr ),
       .io_deq_bits_tag( mem_cmd_q_io_deq_bits_tag ),
       .io_deq_bits_rw( mem_cmd_q_io_deq_bits_rw )
       //.io_count(  )
  );
  Queue_4 mem_data_q(.clk(clk), .reset(reset),
       .io_enq_ready( mem_data_q_io_enq_ready ),
       .io_enq_valid( T32 ),
       .io_enq_bits_data( T0 ),
       .io_deq_ready( io_mem_req_data_ready ),
       .io_deq_valid( mem_data_q_io_deq_valid ),
       .io_deq_bits_data( mem_data_q_io_deq_bits_data )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(T15) begin
      buf_out <= T30;
    end else if(T3) begin
      buf_out <= io_uncached_acquire_bits_payload_data;
    end
    if(reset) begin
      active_out <= 1'h0;
    end else if(T8) begin
      active_out <= 1'h0;
    end else if(T3) begin
      active_out <= 1'h1;
    end
    if(T15) begin
      cnt_out <= T14;
    end else if(T3) begin
      cnt_out <= 3'h0;
    end
    if(reset) begin
      has_data <= 1'h0;
    end else if(T3) begin
      has_data <= T20;
    end
    if(reset) begin
      cmd_sent_out <= 1'h0;
    end else if(T28) begin
      cmd_sent_out <= 1'h1;
    end else if(T3) begin
      cmd_sent_out <= 1'h0;
    end
    if(T3) begin
      tag_out <= io_uncached_acquire_bits_payload_client_xact_id;
    end
    if(T3) begin
      addr_out <= io_uncached_acquire_bits_payload_addr;
    end
    if(T52) begin
      cnt_in <= T51;
    end else if(T44) begin
      cnt_in <= 3'h1;
    end
    if(reset) begin
      active_in <= 1'h0;
    end else if(T49) begin
      active_in <= 1'h0;
    end else if(T44) begin
      active_in <= 1'h1;
    end
    if(T44) begin
      tag_in <= io_mem_resp_bits_tag;
    end
    if(T52) begin
      buf_in <= T64;
    end else if(T44) begin
      buf_in <= T63;
    end
  end
endmodule

module Queue_5(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [4:0] io_enq_bits_tag,
    input  io_enq_bits_rw,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[4:0] io_deq_bits_tag,
    output io_deq_bits_rw
);

  wire T0;
  wire[31:0] T1;
  wire[5:0] T2;
  wire T3;
  wire[31:0] T4;
  reg [31:0] ram [1:0];
  wire[31:0] T5;
  wire[31:0] T6;
  wire[31:0] T7;
  wire[5:0] T8;
  wire do_enq;
  wire T9;
  wire do_flow;
  wire T10;
  reg  enq_ptr;
  wire T11;
  wire T12;
  wire T13;
  reg  deq_ptr;
  wire T14;
  wire T15;
  wire T16;
  wire do_deq;
  wire T17;
  wire T18;
  wire[4:0] T19;
  wire[25:0] T20;
  wire[4:0] T21;
  wire[25:0] T22;
  wire T23;
  wire empty;
  wire T24;
  reg  maybe_full;
  wire T25;
  wire T26;
  wire T27;
  wire ptr_match;
  wire T28;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    enq_ptr = {1{$random}};
    deq_ptr = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_rw = T0;
  assign T0 = T1[1'h0:1'h0];
  assign T1 = {T20, T2};
  assign T2 = {T19, T3};
  assign T3 = T4[1'h0:1'h0];
  assign T4 = ram[deq_ptr];
  always @(posedge clk)
    if (do_enq)
      ram[enq_ptr] <= T6;
  assign T6 = T7;
  assign T7 = {io_enq_bits_addr, T8};
  assign T8 = {io_enq_bits_tag, io_enq_bits_rw};
  assign do_enq = T10 & T9;
  assign T9 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T10 = io_enq_ready & io_enq_valid;
  assign T11 = reset ? 1'h0 : T12;
  assign T12 = do_enq ? T13 : enq_ptr;
  assign T13 = enq_ptr + 1'h1;
  assign T14 = reset ? 1'h0 : T15;
  assign T15 = do_deq ? T16 : deq_ptr;
  assign T16 = deq_ptr + 1'h1;
  assign do_deq = T18 & T17;
  assign T17 = do_flow ^ 1'h1;
  assign T18 = io_deq_ready & io_deq_valid;
  assign T19 = T4[3'h5:1'h1];
  assign T20 = T4[5'h1f:3'h6];
  assign io_deq_bits_tag = T21;
  assign T21 = T1[3'h5:1'h1];
  assign io_deq_bits_addr = T22;
  assign T22 = T1[5'h1f:3'h6];
  assign io_deq_valid = T23;
  assign T23 = empty ^ 1'h1;
  assign empty = ptr_match & T24;
  assign T24 = maybe_full ^ 1'h1;
  assign T25 = reset ? 1'h0 : T26;
  assign T26 = T27 ? do_enq : maybe_full;
  assign T27 = do_enq != do_deq;
  assign ptr_match = enq_ptr == deq_ptr;
  assign io_enq_ready = T28;
  assign T28 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      enq_ptr <= 1'h0;
    end else if(do_enq) begin
      enq_ptr <= T13;
    end
    if(reset) begin
      deq_ptr <= 1'h0;
    end else if(do_deq) begin
      deq_ptr <= T16;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T27) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_6(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data
);

  wire[127:0] T0;
  wire[127:0] T1;
  reg [127:0] ram [3:0];
  wire[127:0] T2;
  wire do_enq;
  wire T3;
  wire do_flow;
  wire T4;
  reg [1:0] enq_ptr;
  wire[1:0] T5;
  wire[1:0] T6;
  wire[1:0] T7;
  reg [1:0] deq_ptr;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire do_deq;
  wire T11;
  wire T12;
  wire T13;
  wire empty;
  wire T14;
  reg  maybe_full;
  wire T15;
  wire T16;
  wire T17;
  wire ptr_match;
  wire T18;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      ram[initvar] = {4{$random}};
    enq_ptr = {1{$random}};
    deq_ptr = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_data = T0;
  assign T0 = T1[7'h7f:1'h0];
  assign T1 = ram[deq_ptr];
  always @(posedge clk)
    if (do_enq)
      ram[enq_ptr] <= io_enq_bits_data;
  assign do_enq = T4 & T3;
  assign T3 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T4 = io_enq_ready & io_enq_valid;
  assign T5 = reset ? 2'h0 : T6;
  assign T6 = do_enq ? T7 : enq_ptr;
  assign T7 = enq_ptr + 2'h1;
  assign T8 = reset ? 2'h0 : T9;
  assign T9 = do_deq ? T10 : deq_ptr;
  assign T10 = deq_ptr + 2'h1;
  assign do_deq = T12 & T11;
  assign T11 = do_flow ^ 1'h1;
  assign T12 = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T13;
  assign T13 = empty ^ 1'h1;
  assign empty = ptr_match & T14;
  assign T14 = maybe_full ^ 1'h1;
  assign T15 = reset ? 1'h0 : T16;
  assign T16 = T17 ? do_enq : maybe_full;
  assign T17 = do_enq != do_deq;
  assign ptr_match = enq_ptr == deq_ptr;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      enq_ptr <= 2'h0;
    end else if(do_enq) begin
      enq_ptr <= T7;
    end
    if(reset) begin
      deq_ptr <= 2'h0;
    end else if(do_deq) begin
      deq_ptr <= T10;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T17) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_7(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input [4:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[4:0] io_deq_bits_tag
);

  wire[4:0] T0;
  wire[132:0] T1;
  wire[4:0] T2;
  wire[132:0] T3;
  reg [132:0] ram [1:0];
  wire[132:0] T4;
  wire[132:0] T5;
  wire[132:0] T6;
  wire do_enq;
  wire T7;
  wire do_flow;
  wire T8;
  reg  enq_ptr;
  wire T9;
  wire T10;
  wire T11;
  reg  deq_ptr;
  wire T12;
  wire T13;
  wire T14;
  wire do_deq;
  wire T15;
  wire T16;
  wire[127:0] T17;
  wire[127:0] T18;
  wire T19;
  wire empty;
  wire T20;
  reg  maybe_full;
  wire T21;
  wire T22;
  wire T23;
  wire ptr_match;
  wire T24;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {5{$random}};
    enq_ptr = {1{$random}};
    deq_ptr = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_tag = T0;
  assign T0 = T1[3'h4:1'h0];
  assign T1 = {T17, T2};
  assign T2 = T3[3'h4:1'h0];
  assign T3 = ram[deq_ptr];
  always @(posedge clk)
    if (do_enq)
      ram[enq_ptr] <= T5;
  assign T5 = T6;
  assign T6 = {io_enq_bits_data, io_enq_bits_tag};
  assign do_enq = T8 & T7;
  assign T7 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T8 = io_enq_ready & io_enq_valid;
  assign T9 = reset ? 1'h0 : T10;
  assign T10 = do_enq ? T11 : enq_ptr;
  assign T11 = enq_ptr + 1'h1;
  assign T12 = reset ? 1'h0 : T13;
  assign T13 = do_deq ? T14 : deq_ptr;
  assign T14 = deq_ptr + 1'h1;
  assign do_deq = T16 & T15;
  assign T15 = do_flow ^ 1'h1;
  assign T16 = io_deq_ready & io_deq_valid;
  assign T17 = T3[8'h84:3'h5];
  assign io_deq_bits_data = T18;
  assign T18 = T1[8'h84:3'h5];
  assign io_deq_valid = T19;
  assign T19 = empty ^ 1'h1;
  assign empty = ptr_match & T20;
  assign T20 = maybe_full ^ 1'h1;
  assign T21 = reset ? 1'h0 : T22;
  assign T22 = T23 ? do_enq : maybe_full;
  assign T23 = do_enq != do_deq;
  assign ptr_match = enq_ptr == deq_ptr;
  assign io_enq_ready = T24;
  assign T24 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      enq_ptr <= 1'h0;
    end else if(do_enq) begin
      enq_ptr <= T11;
    end
    if(reset) begin
      deq_ptr <= 1'h0;
    end else if(do_deq) begin
      deq_ptr <= T14;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T23) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module FPGAOuterMemorySystem(input clk, input reset,
    output io_tiles_0_acquire_ready,
    input  io_tiles_0_acquire_valid,
    input [1:0] io_tiles_0_acquire_bits_header_src,
    input [1:0] io_tiles_0_acquire_bits_header_dst,
    input [25:0] io_tiles_0_acquire_bits_payload_addr,
    input [3:0] io_tiles_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_tiles_0_acquire_bits_payload_data,
    input [2:0] io_tiles_0_acquire_bits_payload_a_type,
    input [5:0] io_tiles_0_acquire_bits_payload_write_mask,
    input [2:0] io_tiles_0_acquire_bits_payload_subword_addr,
    input [3:0] io_tiles_0_acquire_bits_payload_atomic_opcode,
    input  io_tiles_0_grant_ready,
    output io_tiles_0_grant_valid,
    output[1:0] io_tiles_0_grant_bits_header_src,
    output[1:0] io_tiles_0_grant_bits_header_dst,
    output[511:0] io_tiles_0_grant_bits_payload_data,
    output[3:0] io_tiles_0_grant_bits_payload_client_xact_id,
    output[3:0] io_tiles_0_grant_bits_payload_master_xact_id,
    output[3:0] io_tiles_0_grant_bits_payload_g_type,
    output io_tiles_0_finish_ready,
    input  io_tiles_0_finish_valid,
    input [1:0] io_tiles_0_finish_bits_header_src,
    input [1:0] io_tiles_0_finish_bits_header_dst,
    input [3:0] io_tiles_0_finish_bits_payload_master_xact_id,
    input  io_tiles_0_probe_ready,
    output io_tiles_0_probe_valid,
    output[1:0] io_tiles_0_probe_bits_header_src,
    output[1:0] io_tiles_0_probe_bits_header_dst,
    output[25:0] io_tiles_0_probe_bits_payload_addr,
    output[3:0] io_tiles_0_probe_bits_payload_master_xact_id,
    output[1:0] io_tiles_0_probe_bits_payload_p_type,
    output io_tiles_0_release_ready,
    input  io_tiles_0_release_valid,
    input [1:0] io_tiles_0_release_bits_header_src,
    input [1:0] io_tiles_0_release_bits_header_dst,
    input [25:0] io_tiles_0_release_bits_payload_addr,
    input [3:0] io_tiles_0_release_bits_payload_client_xact_id,
    input [3:0] io_tiles_0_release_bits_payload_master_xact_id,
    input [511:0] io_tiles_0_release_bits_payload_data,
    input [2:0] io_tiles_0_release_bits_payload_r_type,
    output io_htif_acquire_ready,
    input  io_htif_acquire_valid,
    input [1:0] io_htif_acquire_bits_header_src,
    input [1:0] io_htif_acquire_bits_header_dst,
    input [25:0] io_htif_acquire_bits_payload_addr,
    input [3:0] io_htif_acquire_bits_payload_client_xact_id,
    input [511:0] io_htif_acquire_bits_payload_data,
    input [2:0] io_htif_acquire_bits_payload_a_type,
    input [5:0] io_htif_acquire_bits_payload_write_mask,
    input [2:0] io_htif_acquire_bits_payload_subword_addr,
    input [3:0] io_htif_acquire_bits_payload_atomic_opcode,
    input  io_htif_grant_ready,
    output io_htif_grant_valid,
    output[1:0] io_htif_grant_bits_header_src,
    output[1:0] io_htif_grant_bits_header_dst,
    output[511:0] io_htif_grant_bits_payload_data,
    output[3:0] io_htif_grant_bits_payload_client_xact_id,
    output[3:0] io_htif_grant_bits_payload_master_xact_id,
    output[3:0] io_htif_grant_bits_payload_g_type,
    output io_htif_finish_ready,
    input  io_htif_finish_valid,
    input [1:0] io_htif_finish_bits_header_src,
    input [1:0] io_htif_finish_bits_header_dst,
    input [3:0] io_htif_finish_bits_payload_master_xact_id,
    input  io_htif_probe_ready,
    output io_htif_probe_valid,
    output[1:0] io_htif_probe_bits_header_src,
    output[1:0] io_htif_probe_bits_header_dst,
    output[25:0] io_htif_probe_bits_payload_addr,
    output[3:0] io_htif_probe_bits_payload_master_xact_id,
    output[1:0] io_htif_probe_bits_payload_p_type,
    output io_htif_release_ready,
    input  io_htif_release_valid,
    input [1:0] io_htif_release_bits_header_src,
    input [1:0] io_htif_release_bits_header_dst,
    input [25:0] io_htif_release_bits_payload_addr,
    input [3:0] io_htif_release_bits_payload_client_xact_id,
    input [3:0] io_htif_release_bits_payload_master_xact_id,
    input [511:0] io_htif_release_bits_payload_data,
    input [2:0] io_htif_release_bits_payload_r_type,
    input  io_incoherent_1,
    input  io_incoherent_0,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    output io_mem_resp_ready,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
);

  wire conv_io_mem_resp_ready;
  wire[127:0] conv_io_mem_req_data_bits_data;
  wire conv_io_mem_req_data_valid;
  wire conv_io_mem_req_cmd_bits_rw;
  wire[4:0] conv_io_mem_req_cmd_bits_tag;
  wire[25:0] conv_io_mem_req_cmd_bits_addr;
  wire conv_io_mem_req_cmd_valid;
  wire[4:0] Queue_2_io_deq_bits_tag;
  wire[127:0] Queue_2_io_deq_bits_data;
  wire Queue_2_io_deq_valid;
  wire Queue_1_io_enq_ready;
  wire Queue_0_io_enq_ready;
  wire[3:0] master_io_outer_finish_bits_payload_master_xact_id;
  wire[1:0] master_io_outer_finish_bits_header_dst;
  wire[1:0] master_io_outer_finish_bits_header_src;
  wire master_io_outer_finish_valid;
  wire master_io_outer_grant_ready;
  wire[3:0] master_io_outer_acquire_bits_payload_atomic_opcode;
  wire[2:0] master_io_outer_acquire_bits_payload_subword_addr;
  wire[5:0] master_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] master_io_outer_acquire_bits_payload_a_type;
  wire[511:0] master_io_outer_acquire_bits_payload_data;
  wire[3:0] master_io_outer_acquire_bits_payload_client_xact_id;
  wire[25:0] master_io_outer_acquire_bits_payload_addr;
  wire[1:0] master_io_outer_acquire_bits_header_dst;
  wire[1:0] master_io_outer_acquire_bits_header_src;
  wire master_io_outer_acquire_valid;
  wire master_io_inner_release_ready;
  wire[1:0] master_io_inner_probe_bits_payload_p_type;
  wire[3:0] master_io_inner_probe_bits_payload_master_xact_id;
  wire[25:0] master_io_inner_probe_bits_payload_addr;
  wire[1:0] master_io_inner_probe_bits_header_dst;
  wire[1:0] master_io_inner_probe_bits_header_src;
  wire master_io_inner_probe_valid;
  wire master_io_inner_finish_ready;
  wire[3:0] master_io_inner_grant_bits_payload_g_type;
  wire[3:0] master_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] master_io_inner_grant_bits_payload_client_xact_id;
  wire[511:0] master_io_inner_grant_bits_payload_data;
  wire[1:0] master_io_inner_grant_bits_header_dst;
  wire[1:0] master_io_inner_grant_bits_header_src;
  wire master_io_inner_grant_valid;
  wire master_io_inner_acquire_ready;
  wire[3:0] conv_io_uncached_grant_bits_payload_g_type;
  wire[3:0] conv_io_uncached_grant_bits_payload_master_xact_id;
  wire[3:0] conv_io_uncached_grant_bits_payload_client_xact_id;
  wire[511:0] conv_io_uncached_grant_bits_payload_data;
  wire conv_io_uncached_grant_valid;
  wire conv_io_uncached_acquire_ready;
  wire[2:0] net_io_masters_0_release_bits_payload_r_type;
  wire[511:0] net_io_masters_0_release_bits_payload_data;
  wire[3:0] net_io_masters_0_release_bits_payload_master_xact_id;
  wire[3:0] net_io_masters_0_release_bits_payload_client_xact_id;
  wire[25:0] net_io_masters_0_release_bits_payload_addr;
  wire[1:0] net_io_masters_0_release_bits_header_dst;
  wire[1:0] net_io_masters_0_release_bits_header_src;
  wire net_io_masters_0_release_valid;
  wire net_io_masters_0_probe_ready;
  wire[3:0] net_io_masters_0_finish_bits_payload_master_xact_id;
  wire[1:0] net_io_masters_0_finish_bits_header_dst;
  wire[1:0] net_io_masters_0_finish_bits_header_src;
  wire net_io_masters_0_finish_valid;
  wire net_io_masters_0_grant_ready;
  wire[3:0] net_io_masters_0_acquire_bits_payload_atomic_opcode;
  wire[2:0] net_io_masters_0_acquire_bits_payload_subword_addr;
  wire[5:0] net_io_masters_0_acquire_bits_payload_write_mask;
  wire[2:0] net_io_masters_0_acquire_bits_payload_a_type;
  wire[511:0] net_io_masters_0_acquire_bits_payload_data;
  wire[3:0] net_io_masters_0_acquire_bits_payload_client_xact_id;
  wire[25:0] net_io_masters_0_acquire_bits_payload_addr;
  wire[1:0] net_io_masters_0_acquire_bits_header_dst;
  wire[1:0] net_io_masters_0_acquire_bits_header_src;
  wire net_io_masters_0_acquire_valid;
  wire Queue_2_io_enq_ready;
  wire[127:0] Queue_1_io_deq_bits_data;
  wire Queue_1_io_deq_valid;
  wire Queue_0_io_deq_bits_rw;
  wire[4:0] Queue_0_io_deq_bits_tag;
  wire[25:0] Queue_0_io_deq_bits_addr;
  wire Queue_0_io_deq_valid;
  wire net_io_clients_1_release_ready;
  wire[1:0] net_io_clients_1_probe_bits_payload_p_type;
  wire[3:0] net_io_clients_1_probe_bits_payload_master_xact_id;
  wire[25:0] net_io_clients_1_probe_bits_payload_addr;
  wire[1:0] net_io_clients_1_probe_bits_header_dst;
  wire[1:0] net_io_clients_1_probe_bits_header_src;
  wire net_io_clients_1_probe_valid;
  wire net_io_clients_1_finish_ready;
  wire[3:0] net_io_clients_1_grant_bits_payload_g_type;
  wire[3:0] net_io_clients_1_grant_bits_payload_master_xact_id;
  wire[3:0] net_io_clients_1_grant_bits_payload_client_xact_id;
  wire[511:0] net_io_clients_1_grant_bits_payload_data;
  wire[1:0] net_io_clients_1_grant_bits_header_dst;
  wire[1:0] net_io_clients_1_grant_bits_header_src;
  wire net_io_clients_1_grant_valid;
  wire net_io_clients_1_acquire_ready;
  wire net_io_clients_0_release_ready;
  wire[1:0] net_io_clients_0_probe_bits_payload_p_type;
  wire[3:0] net_io_clients_0_probe_bits_payload_master_xact_id;
  wire[25:0] net_io_clients_0_probe_bits_payload_addr;
  wire[1:0] net_io_clients_0_probe_bits_header_dst;
  wire[1:0] net_io_clients_0_probe_bits_header_src;
  wire net_io_clients_0_probe_valid;
  wire net_io_clients_0_finish_ready;
  wire[3:0] net_io_clients_0_grant_bits_payload_g_type;
  wire[3:0] net_io_clients_0_grant_bits_payload_master_xact_id;
  wire[3:0] net_io_clients_0_grant_bits_payload_client_xact_id;
  wire[511:0] net_io_clients_0_grant_bits_payload_data;
  wire[1:0] net_io_clients_0_grant_bits_header_dst;
  wire[1:0] net_io_clients_0_grant_bits_header_src;
  wire net_io_clients_0_grant_valid;
  wire net_io_clients_0_acquire_ready;


  assign io_mem_resp_ready = Queue_2_io_enq_ready;
  assign io_mem_req_data_bits_data = Queue_1_io_deq_bits_data;
  assign io_mem_req_data_valid = Queue_1_io_deq_valid;
  assign io_mem_req_cmd_bits_rw = Queue_0_io_deq_bits_rw;
  assign io_mem_req_cmd_bits_tag = Queue_0_io_deq_bits_tag;
  assign io_mem_req_cmd_bits_addr = Queue_0_io_deq_bits_addr;
  assign io_mem_req_cmd_valid = Queue_0_io_deq_valid;
  assign io_htif_release_ready = net_io_clients_1_release_ready;
  assign io_htif_probe_bits_payload_p_type = net_io_clients_1_probe_bits_payload_p_type;
  assign io_htif_probe_bits_payload_master_xact_id = net_io_clients_1_probe_bits_payload_master_xact_id;
  assign io_htif_probe_bits_payload_addr = net_io_clients_1_probe_bits_payload_addr;
  assign io_htif_probe_bits_header_dst = net_io_clients_1_probe_bits_header_dst;
  assign io_htif_probe_bits_header_src = net_io_clients_1_probe_bits_header_src;
  assign io_htif_probe_valid = net_io_clients_1_probe_valid;
  assign io_htif_finish_ready = net_io_clients_1_finish_ready;
  assign io_htif_grant_bits_payload_g_type = net_io_clients_1_grant_bits_payload_g_type;
  assign io_htif_grant_bits_payload_master_xact_id = net_io_clients_1_grant_bits_payload_master_xact_id;
  assign io_htif_grant_bits_payload_client_xact_id = net_io_clients_1_grant_bits_payload_client_xact_id;
  assign io_htif_grant_bits_payload_data = net_io_clients_1_grant_bits_payload_data;
  assign io_htif_grant_bits_header_dst = net_io_clients_1_grant_bits_header_dst;
  assign io_htif_grant_bits_header_src = net_io_clients_1_grant_bits_header_src;
  assign io_htif_grant_valid = net_io_clients_1_grant_valid;
  assign io_htif_acquire_ready = net_io_clients_1_acquire_ready;
  assign io_tiles_0_release_ready = net_io_clients_0_release_ready;
  assign io_tiles_0_probe_bits_payload_p_type = net_io_clients_0_probe_bits_payload_p_type;
  assign io_tiles_0_probe_bits_payload_master_xact_id = net_io_clients_0_probe_bits_payload_master_xact_id;
  assign io_tiles_0_probe_bits_payload_addr = net_io_clients_0_probe_bits_payload_addr;
  assign io_tiles_0_probe_bits_header_dst = net_io_clients_0_probe_bits_header_dst;
  assign io_tiles_0_probe_bits_header_src = net_io_clients_0_probe_bits_header_src;
  assign io_tiles_0_probe_valid = net_io_clients_0_probe_valid;
  assign io_tiles_0_finish_ready = net_io_clients_0_finish_ready;
  assign io_tiles_0_grant_bits_payload_g_type = net_io_clients_0_grant_bits_payload_g_type;
  assign io_tiles_0_grant_bits_payload_master_xact_id = net_io_clients_0_grant_bits_payload_master_xact_id;
  assign io_tiles_0_grant_bits_payload_client_xact_id = net_io_clients_0_grant_bits_payload_client_xact_id;
  assign io_tiles_0_grant_bits_payload_data = net_io_clients_0_grant_bits_payload_data;
  assign io_tiles_0_grant_bits_header_dst = net_io_clients_0_grant_bits_header_dst;
  assign io_tiles_0_grant_bits_header_src = net_io_clients_0_grant_bits_header_src;
  assign io_tiles_0_grant_valid = net_io_clients_0_grant_valid;
  assign io_tiles_0_acquire_ready = net_io_clients_0_acquire_ready;
  L2CoherenceAgent master(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( master_io_inner_acquire_ready ),
       .io_inner_acquire_valid( net_io_masters_0_acquire_valid ),
       .io_inner_acquire_bits_header_src( net_io_masters_0_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( net_io_masters_0_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( net_io_masters_0_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( net_io_masters_0_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( net_io_masters_0_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( net_io_masters_0_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( net_io_masters_0_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( net_io_masters_0_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( net_io_masters_0_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( net_io_masters_0_grant_ready ),
       .io_inner_grant_valid( master_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( master_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( master_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( master_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( master_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( master_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( master_io_inner_grant_bits_payload_g_type ),
       .io_inner_finish_ready( master_io_inner_finish_ready ),
       .io_inner_finish_valid( net_io_masters_0_finish_valid ),
       .io_inner_finish_bits_header_src( net_io_masters_0_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( net_io_masters_0_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( net_io_masters_0_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( net_io_masters_0_probe_ready ),
       .io_inner_probe_valid( master_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( master_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( master_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( master_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( master_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( master_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( master_io_inner_release_ready ),
       .io_inner_release_valid( net_io_masters_0_release_valid ),
       .io_inner_release_bits_header_src( net_io_masters_0_release_bits_header_src ),
       .io_inner_release_bits_header_dst( net_io_masters_0_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( net_io_masters_0_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( net_io_masters_0_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( net_io_masters_0_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( net_io_masters_0_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( net_io_masters_0_release_bits_payload_r_type ),
       .io_outer_acquire_ready( conv_io_uncached_acquire_ready ),
       .io_outer_acquire_valid( master_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( master_io_outer_acquire_bits_header_src ),
       .io_outer_acquire_bits_header_dst( master_io_outer_acquire_bits_header_dst ),
       .io_outer_acquire_bits_payload_addr( master_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( master_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( master_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( master_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( master_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( master_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( master_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( master_io_outer_grant_ready ),
       .io_outer_grant_valid( conv_io_uncached_grant_valid ),
       //.io_outer_grant_bits_header_src(  )
       //.io_outer_grant_bits_header_dst(  )
       .io_outer_grant_bits_payload_data( conv_io_uncached_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( conv_io_uncached_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( conv_io_uncached_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( conv_io_uncached_grant_bits_payload_g_type ),
       //.io_outer_finish_ready(  )
       .io_outer_finish_valid( master_io_outer_finish_valid ),
       .io_outer_finish_bits_header_src( master_io_outer_finish_bits_header_src ),
       .io_outer_finish_bits_header_dst( master_io_outer_finish_bits_header_dst ),
       .io_outer_finish_bits_payload_master_xact_id( master_io_outer_finish_bits_payload_master_xact_id ),
       .io_incoherent_1( io_incoherent_1 ),
       .io_incoherent_0( io_incoherent_0 )
  );
  `ifndef SYNTHESIS
    assign master.io_outer_grant_bits_header_src = {1{$random}};
    assign master.io_outer_grant_bits_header_dst = {1{$random}};
    assign master.io_outer_finish_ready = {1{$random}};
  `endif
  ReferenceChipCrossbarNetwork net(.clk(clk), .reset(reset),
       .io_clients_1_acquire_ready( net_io_clients_1_acquire_ready ),
       .io_clients_1_acquire_valid( io_htif_acquire_valid ),
       .io_clients_1_acquire_bits_header_src( io_htif_acquire_bits_header_src ),
       .io_clients_1_acquire_bits_header_dst( io_htif_acquire_bits_header_dst ),
       .io_clients_1_acquire_bits_payload_addr( io_htif_acquire_bits_payload_addr ),
       .io_clients_1_acquire_bits_payload_client_xact_id( io_htif_acquire_bits_payload_client_xact_id ),
       .io_clients_1_acquire_bits_payload_data( io_htif_acquire_bits_payload_data ),
       .io_clients_1_acquire_bits_payload_a_type( io_htif_acquire_bits_payload_a_type ),
       .io_clients_1_acquire_bits_payload_write_mask( io_htif_acquire_bits_payload_write_mask ),
       .io_clients_1_acquire_bits_payload_subword_addr( io_htif_acquire_bits_payload_subword_addr ),
       .io_clients_1_acquire_bits_payload_atomic_opcode( io_htif_acquire_bits_payload_atomic_opcode ),
       .io_clients_1_grant_ready( io_htif_grant_ready ),
       .io_clients_1_grant_valid( net_io_clients_1_grant_valid ),
       .io_clients_1_grant_bits_header_src( net_io_clients_1_grant_bits_header_src ),
       .io_clients_1_grant_bits_header_dst( net_io_clients_1_grant_bits_header_dst ),
       .io_clients_1_grant_bits_payload_data( net_io_clients_1_grant_bits_payload_data ),
       .io_clients_1_grant_bits_payload_client_xact_id( net_io_clients_1_grant_bits_payload_client_xact_id ),
       .io_clients_1_grant_bits_payload_master_xact_id( net_io_clients_1_grant_bits_payload_master_xact_id ),
       .io_clients_1_grant_bits_payload_g_type( net_io_clients_1_grant_bits_payload_g_type ),
       .io_clients_1_finish_ready( net_io_clients_1_finish_ready ),
       .io_clients_1_finish_valid( io_htif_finish_valid ),
       .io_clients_1_finish_bits_header_src( io_htif_finish_bits_header_src ),
       .io_clients_1_finish_bits_header_dst( io_htif_finish_bits_header_dst ),
       .io_clients_1_finish_bits_payload_master_xact_id( io_htif_finish_bits_payload_master_xact_id ),
       .io_clients_1_probe_ready( io_htif_probe_ready ),
       .io_clients_1_probe_valid( net_io_clients_1_probe_valid ),
       .io_clients_1_probe_bits_header_src( net_io_clients_1_probe_bits_header_src ),
       .io_clients_1_probe_bits_header_dst( net_io_clients_1_probe_bits_header_dst ),
       .io_clients_1_probe_bits_payload_addr( net_io_clients_1_probe_bits_payload_addr ),
       .io_clients_1_probe_bits_payload_master_xact_id( net_io_clients_1_probe_bits_payload_master_xact_id ),
       .io_clients_1_probe_bits_payload_p_type( net_io_clients_1_probe_bits_payload_p_type ),
       .io_clients_1_release_ready( net_io_clients_1_release_ready ),
       .io_clients_1_release_valid( io_htif_release_valid ),
       .io_clients_1_release_bits_header_src( io_htif_release_bits_header_src ),
       .io_clients_1_release_bits_header_dst( io_htif_release_bits_header_dst ),
       .io_clients_1_release_bits_payload_addr( io_htif_release_bits_payload_addr ),
       .io_clients_1_release_bits_payload_client_xact_id( io_htif_release_bits_payload_client_xact_id ),
       .io_clients_1_release_bits_payload_master_xact_id( io_htif_release_bits_payload_master_xact_id ),
       .io_clients_1_release_bits_payload_data( io_htif_release_bits_payload_data ),
       .io_clients_1_release_bits_payload_r_type( io_htif_release_bits_payload_r_type ),
       .io_clients_0_acquire_ready( net_io_clients_0_acquire_ready ),
       .io_clients_0_acquire_valid( io_tiles_0_acquire_valid ),
       .io_clients_0_acquire_bits_header_src( io_tiles_0_acquire_bits_header_src ),
       .io_clients_0_acquire_bits_header_dst( io_tiles_0_acquire_bits_header_dst ),
       .io_clients_0_acquire_bits_payload_addr( io_tiles_0_acquire_bits_payload_addr ),
       .io_clients_0_acquire_bits_payload_client_xact_id( io_tiles_0_acquire_bits_payload_client_xact_id ),
       .io_clients_0_acquire_bits_payload_data( io_tiles_0_acquire_bits_payload_data ),
       .io_clients_0_acquire_bits_payload_a_type( io_tiles_0_acquire_bits_payload_a_type ),
       .io_clients_0_acquire_bits_payload_write_mask( io_tiles_0_acquire_bits_payload_write_mask ),
       .io_clients_0_acquire_bits_payload_subword_addr( io_tiles_0_acquire_bits_payload_subword_addr ),
       .io_clients_0_acquire_bits_payload_atomic_opcode( io_tiles_0_acquire_bits_payload_atomic_opcode ),
       .io_clients_0_grant_ready( io_tiles_0_grant_ready ),
       .io_clients_0_grant_valid( net_io_clients_0_grant_valid ),
       .io_clients_0_grant_bits_header_src( net_io_clients_0_grant_bits_header_src ),
       .io_clients_0_grant_bits_header_dst( net_io_clients_0_grant_bits_header_dst ),
       .io_clients_0_grant_bits_payload_data( net_io_clients_0_grant_bits_payload_data ),
       .io_clients_0_grant_bits_payload_client_xact_id( net_io_clients_0_grant_bits_payload_client_xact_id ),
       .io_clients_0_grant_bits_payload_master_xact_id( net_io_clients_0_grant_bits_payload_master_xact_id ),
       .io_clients_0_grant_bits_payload_g_type( net_io_clients_0_grant_bits_payload_g_type ),
       .io_clients_0_finish_ready( net_io_clients_0_finish_ready ),
       .io_clients_0_finish_valid( io_tiles_0_finish_valid ),
       .io_clients_0_finish_bits_header_src( io_tiles_0_finish_bits_header_src ),
       .io_clients_0_finish_bits_header_dst( io_tiles_0_finish_bits_header_dst ),
       .io_clients_0_finish_bits_payload_master_xact_id( io_tiles_0_finish_bits_payload_master_xact_id ),
       .io_clients_0_probe_ready( io_tiles_0_probe_ready ),
       .io_clients_0_probe_valid( net_io_clients_0_probe_valid ),
       .io_clients_0_probe_bits_header_src( net_io_clients_0_probe_bits_header_src ),
       .io_clients_0_probe_bits_header_dst( net_io_clients_0_probe_bits_header_dst ),
       .io_clients_0_probe_bits_payload_addr( net_io_clients_0_probe_bits_payload_addr ),
       .io_clients_0_probe_bits_payload_master_xact_id( net_io_clients_0_probe_bits_payload_master_xact_id ),
       .io_clients_0_probe_bits_payload_p_type( net_io_clients_0_probe_bits_payload_p_type ),
       .io_clients_0_release_ready( net_io_clients_0_release_ready ),
       .io_clients_0_release_valid( io_tiles_0_release_valid ),
       .io_clients_0_release_bits_header_src( io_tiles_0_release_bits_header_src ),
       .io_clients_0_release_bits_header_dst( io_tiles_0_release_bits_header_dst ),
       .io_clients_0_release_bits_payload_addr( io_tiles_0_release_bits_payload_addr ),
       .io_clients_0_release_bits_payload_client_xact_id( io_tiles_0_release_bits_payload_client_xact_id ),
       .io_clients_0_release_bits_payload_master_xact_id( io_tiles_0_release_bits_payload_master_xact_id ),
       .io_clients_0_release_bits_payload_data( io_tiles_0_release_bits_payload_data ),
       .io_clients_0_release_bits_payload_r_type( io_tiles_0_release_bits_payload_r_type ),
       .io_masters_0_acquire_ready( master_io_inner_acquire_ready ),
       .io_masters_0_acquire_valid( net_io_masters_0_acquire_valid ),
       .io_masters_0_acquire_bits_header_src( net_io_masters_0_acquire_bits_header_src ),
       .io_masters_0_acquire_bits_header_dst( net_io_masters_0_acquire_bits_header_dst ),
       .io_masters_0_acquire_bits_payload_addr( net_io_masters_0_acquire_bits_payload_addr ),
       .io_masters_0_acquire_bits_payload_client_xact_id( net_io_masters_0_acquire_bits_payload_client_xact_id ),
       .io_masters_0_acquire_bits_payload_data( net_io_masters_0_acquire_bits_payload_data ),
       .io_masters_0_acquire_bits_payload_a_type( net_io_masters_0_acquire_bits_payload_a_type ),
       .io_masters_0_acquire_bits_payload_write_mask( net_io_masters_0_acquire_bits_payload_write_mask ),
       .io_masters_0_acquire_bits_payload_subword_addr( net_io_masters_0_acquire_bits_payload_subword_addr ),
       .io_masters_0_acquire_bits_payload_atomic_opcode( net_io_masters_0_acquire_bits_payload_atomic_opcode ),
       .io_masters_0_grant_ready( net_io_masters_0_grant_ready ),
       .io_masters_0_grant_valid( master_io_inner_grant_valid ),
       .io_masters_0_grant_bits_header_src( master_io_inner_grant_bits_header_src ),
       .io_masters_0_grant_bits_header_dst( master_io_inner_grant_bits_header_dst ),
       .io_masters_0_grant_bits_payload_data( master_io_inner_grant_bits_payload_data ),
       .io_masters_0_grant_bits_payload_client_xact_id( master_io_inner_grant_bits_payload_client_xact_id ),
       .io_masters_0_grant_bits_payload_master_xact_id( master_io_inner_grant_bits_payload_master_xact_id ),
       .io_masters_0_grant_bits_payload_g_type( master_io_inner_grant_bits_payload_g_type ),
       .io_masters_0_finish_ready( master_io_inner_finish_ready ),
       .io_masters_0_finish_valid( net_io_masters_0_finish_valid ),
       .io_masters_0_finish_bits_header_src( net_io_masters_0_finish_bits_header_src ),
       .io_masters_0_finish_bits_header_dst( net_io_masters_0_finish_bits_header_dst ),
       .io_masters_0_finish_bits_payload_master_xact_id( net_io_masters_0_finish_bits_payload_master_xact_id ),
       .io_masters_0_probe_ready( net_io_masters_0_probe_ready ),
       .io_masters_0_probe_valid( master_io_inner_probe_valid ),
       .io_masters_0_probe_bits_header_src( master_io_inner_probe_bits_header_src ),
       .io_masters_0_probe_bits_header_dst( master_io_inner_probe_bits_header_dst ),
       .io_masters_0_probe_bits_payload_addr( master_io_inner_probe_bits_payload_addr ),
       .io_masters_0_probe_bits_payload_master_xact_id( master_io_inner_probe_bits_payload_master_xact_id ),
       .io_masters_0_probe_bits_payload_p_type( master_io_inner_probe_bits_payload_p_type ),
       .io_masters_0_release_ready( master_io_inner_release_ready ),
       .io_masters_0_release_valid( net_io_masters_0_release_valid ),
       .io_masters_0_release_bits_header_src( net_io_masters_0_release_bits_header_src ),
       .io_masters_0_release_bits_header_dst( net_io_masters_0_release_bits_header_dst ),
       .io_masters_0_release_bits_payload_addr( net_io_masters_0_release_bits_payload_addr ),
       .io_masters_0_release_bits_payload_client_xact_id( net_io_masters_0_release_bits_payload_client_xact_id ),
       .io_masters_0_release_bits_payload_master_xact_id( net_io_masters_0_release_bits_payload_master_xact_id ),
       .io_masters_0_release_bits_payload_data( net_io_masters_0_release_bits_payload_data ),
       .io_masters_0_release_bits_payload_r_type( net_io_masters_0_release_bits_payload_r_type )
  );
  MemIOUncachedTileLinkIOConverter conv(.clk(clk), .reset(reset),
       .io_uncached_acquire_ready( conv_io_uncached_acquire_ready ),
       .io_uncached_acquire_valid( master_io_outer_acquire_valid ),
       .io_uncached_acquire_bits_header_src( master_io_outer_acquire_bits_header_src ),
       .io_uncached_acquire_bits_header_dst( master_io_outer_acquire_bits_header_dst ),
       .io_uncached_acquire_bits_payload_addr( master_io_outer_acquire_bits_payload_addr ),
       .io_uncached_acquire_bits_payload_client_xact_id( master_io_outer_acquire_bits_payload_client_xact_id ),
       .io_uncached_acquire_bits_payload_data( master_io_outer_acquire_bits_payload_data ),
       .io_uncached_acquire_bits_payload_a_type( master_io_outer_acquire_bits_payload_a_type ),
       .io_uncached_acquire_bits_payload_write_mask( master_io_outer_acquire_bits_payload_write_mask ),
       .io_uncached_acquire_bits_payload_subword_addr( master_io_outer_acquire_bits_payload_subword_addr ),
       .io_uncached_acquire_bits_payload_atomic_opcode( master_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_uncached_grant_ready( master_io_outer_grant_ready ),
       .io_uncached_grant_valid( conv_io_uncached_grant_valid ),
       //.io_uncached_grant_bits_header_src(  )
       //.io_uncached_grant_bits_header_dst(  )
       .io_uncached_grant_bits_payload_data( conv_io_uncached_grant_bits_payload_data ),
       .io_uncached_grant_bits_payload_client_xact_id( conv_io_uncached_grant_bits_payload_client_xact_id ),
       .io_uncached_grant_bits_payload_master_xact_id( conv_io_uncached_grant_bits_payload_master_xact_id ),
       .io_uncached_grant_bits_payload_g_type( conv_io_uncached_grant_bits_payload_g_type ),
       //.io_uncached_finish_ready(  )
       .io_uncached_finish_valid( master_io_outer_finish_valid ),
       .io_uncached_finish_bits_header_src( master_io_outer_finish_bits_header_src ),
       .io_uncached_finish_bits_header_dst( master_io_outer_finish_bits_header_dst ),
       .io_uncached_finish_bits_payload_master_xact_id( master_io_outer_finish_bits_payload_master_xact_id ),
       .io_mem_req_cmd_ready( Queue_0_io_enq_ready ),
       .io_mem_req_cmd_valid( conv_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( conv_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( conv_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( conv_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( Queue_1_io_enq_ready ),
       .io_mem_req_data_valid( conv_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( conv_io_mem_req_data_bits_data ),
       .io_mem_resp_ready( conv_io_mem_resp_ready ),
       .io_mem_resp_valid( Queue_2_io_deq_valid ),
       .io_mem_resp_bits_data( Queue_2_io_deq_bits_data ),
       .io_mem_resp_bits_tag( Queue_2_io_deq_bits_tag )
  );
  Queue_5 Queue_0(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_0_io_enq_ready ),
       .io_enq_valid( conv_io_mem_req_cmd_valid ),
       .io_enq_bits_addr( conv_io_mem_req_cmd_bits_addr ),
       .io_enq_bits_tag( conv_io_mem_req_cmd_bits_tag ),
       .io_enq_bits_rw( conv_io_mem_req_cmd_bits_rw ),
       .io_deq_ready( io_mem_req_cmd_ready ),
       .io_deq_valid( Queue_0_io_deq_valid ),
       .io_deq_bits_addr( Queue_0_io_deq_bits_addr ),
       .io_deq_bits_tag( Queue_0_io_deq_bits_tag ),
       .io_deq_bits_rw( Queue_0_io_deq_bits_rw )
  );
  Queue_6 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( conv_io_mem_req_data_valid ),
       .io_enq_bits_data( conv_io_mem_req_data_bits_data ),
       .io_deq_ready( io_mem_req_data_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits_data( Queue_1_io_deq_bits_data )
  );
  Queue_7 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( io_mem_resp_valid ),
       .io_enq_bits_data( io_mem_resp_bits_data ),
       .io_enq_bits_tag( io_mem_resp_bits_tag ),
       .io_deq_ready( conv_io_mem_resp_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits_data( Queue_2_io_deq_bits_data ),
       .io_deq_bits_tag( Queue_2_io_deq_bits_tag )
  );
endmodule

module Queue_8(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [3:0] io_enq_bits_payload_client_xact_id,
    input [511:0] io_enq_bits_payload_data,
    input [2:0] io_enq_bits_payload_a_type,
    input [5:0] io_enq_bits_payload_write_mask,
    input [2:0] io_enq_bits_payload_subword_addr,
    input [3:0] io_enq_bits_payload_atomic_opcode,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[3:0] io_deq_bits_payload_client_xact_id,
    output[511:0] io_deq_bits_payload_data,
    output[2:0] io_deq_bits_payload_a_type,
    output[5:0] io_deq_bits_payload_write_mask,
    output[2:0] io_deq_bits_payload_subword_addr,
    output[3:0] io_deq_bits_payload_atomic_opcode
);

  wire[3:0] T0;
  wire[561:0] T1;
  wire[527:0] T2;
  wire[12:0] T3;
  wire[6:0] T4;
  wire[3:0] T5;
  wire[561:0] T6;
  reg [561:0] ram [1:0];
  wire[561:0] T7;
  wire[561:0] T8;
  wire[561:0] T9;
  wire[527:0] T10;
  wire[12:0] T11;
  wire[6:0] T12;
  wire[514:0] T13;
  wire[33:0] T14;
  wire[29:0] T15;
  wire[3:0] T16;
  wire do_enq;
  wire T17;
  wire do_flow;
  wire T18;
  reg  enq_ptr;
  wire T19;
  wire T20;
  wire T21;
  reg  deq_ptr;
  wire T22;
  wire T23;
  wire T24;
  wire do_deq;
  wire T25;
  wire T26;
  wire[2:0] T27;
  wire[5:0] T28;
  wire[514:0] T29;
  wire[2:0] T30;
  wire[511:0] T31;
  wire[33:0] T32;
  wire[29:0] T33;
  wire[3:0] T34;
  wire[25:0] T35;
  wire[3:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[2:0] T39;
  wire[5:0] T40;
  wire[2:0] T41;
  wire[511:0] T42;
  wire[3:0] T43;
  wire[25:0] T44;
  wire[1:0] T45;
  wire[1:0] T46;
  wire T47;
  wire empty;
  wire T48;
  reg  maybe_full;
  wire T49;
  wire T50;
  wire T51;
  wire ptr_match;
  wire T52;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {18{$random}};
    enq_ptr = {1{$random}};
    deq_ptr = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_atomic_opcode = T0;
  assign T0 = T1[2'h3:1'h0];
  assign T1 = {T32, T2};
  assign T2 = {T29, T3};
  assign T3 = {T28, T4};
  assign T4 = {T27, T5};
  assign T5 = T6[2'h3:1'h0];
  assign T6 = ram[deq_ptr];
  always @(posedge clk)
    if (do_enq)
      ram[enq_ptr] <= T8;
  assign T8 = T9;
  assign T9 = {T14, T10};
  assign T10 = {T13, T11};
  assign T11 = {io_enq_bits_payload_write_mask, T12};
  assign T12 = {io_enq_bits_payload_subword_addr, io_enq_bits_payload_atomic_opcode};
  assign T13 = {io_enq_bits_payload_data, io_enq_bits_payload_a_type};
  assign T14 = {T16, T15};
  assign T15 = {io_enq_bits_payload_addr, io_enq_bits_payload_client_xact_id};
  assign T16 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign do_enq = T18 & T17;
  assign T17 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T18 = io_enq_ready & io_enq_valid;
  assign T19 = reset ? 1'h0 : T20;
  assign T20 = do_enq ? T21 : enq_ptr;
  assign T21 = enq_ptr + 1'h1;
  assign T22 = reset ? 1'h0 : T23;
  assign T23 = do_deq ? T24 : deq_ptr;
  assign T24 = deq_ptr + 1'h1;
  assign do_deq = T26 & T25;
  assign T25 = do_flow ^ 1'h1;
  assign T26 = io_deq_ready & io_deq_valid;
  assign T27 = T6[3'h6:3'h4];
  assign T28 = T6[4'hc:3'h7];
  assign T29 = {T31, T30};
  assign T30 = T6[4'hf:4'hd];
  assign T31 = T6[10'h20f:5'h10];
  assign T32 = {T36, T33};
  assign T33 = {T35, T34};
  assign T34 = T6[10'h213:10'h210];
  assign T35 = T6[10'h22d:10'h214];
  assign T36 = {T38, T37};
  assign T37 = T6[10'h22f:10'h22e];
  assign T38 = T6[10'h231:10'h230];
  assign io_deq_bits_payload_subword_addr = T39;
  assign T39 = T1[3'h6:3'h4];
  assign io_deq_bits_payload_write_mask = T40;
  assign T40 = T1[4'hc:3'h7];
  assign io_deq_bits_payload_a_type = T41;
  assign T41 = T1[4'hf:4'hd];
  assign io_deq_bits_payload_data = T42;
  assign T42 = T1[10'h20f:5'h10];
  assign io_deq_bits_payload_client_xact_id = T43;
  assign T43 = T1[10'h213:10'h210];
  assign io_deq_bits_payload_addr = T44;
  assign T44 = T1[10'h22d:10'h214];
  assign io_deq_bits_header_dst = T45;
  assign T45 = T1[10'h22f:10'h22e];
  assign io_deq_bits_header_src = T46;
  assign T46 = T1[10'h231:10'h230];
  assign io_deq_valid = T47;
  assign T47 = empty ^ 1'h1;
  assign empty = ptr_match & T48;
  assign T48 = maybe_full ^ 1'h1;
  assign T49 = reset ? 1'h0 : T50;
  assign T50 = T51 ? do_enq : maybe_full;
  assign T51 = do_enq != do_deq;
  assign ptr_match = enq_ptr == deq_ptr;
  assign io_enq_ready = T52;
  assign T52 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      enq_ptr <= 1'h0;
    end else if(do_enq) begin
      enq_ptr <= T21;
    end
    if(reset) begin
      deq_ptr <= 1'h0;
    end else if(do_deq) begin
      deq_ptr <= T24;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T51) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_9(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [3:0] io_enq_bits_payload_client_xact_id,
    input [3:0] io_enq_bits_payload_master_xact_id,
    input [511:0] io_enq_bits_payload_data,
    input [2:0] io_enq_bits_payload_r_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[3:0] io_deq_bits_payload_client_xact_id,
    output[3:0] io_deq_bits_payload_master_xact_id,
    output[511:0] io_deq_bits_payload_data,
    output[2:0] io_deq_bits_payload_r_type
);

  wire[2:0] T0;
  wire[552:0] T1;
  wire[522:0] T2;
  wire[514:0] T3;
  wire[2:0] T4;
  wire[552:0] T5;
  reg [552:0] ram [1:0];
  wire[552:0] T6;
  wire[552:0] T7;
  wire[552:0] T8;
  wire[522:0] T9;
  wire[514:0] T10;
  wire[7:0] T11;
  wire[29:0] T12;
  wire[27:0] T13;
  wire do_enq;
  wire T14;
  wire do_flow;
  wire T15;
  reg  enq_ptr;
  wire T16;
  wire T17;
  wire T18;
  reg  deq_ptr;
  wire T19;
  wire T20;
  wire T21;
  wire do_deq;
  wire T22;
  wire T23;
  wire[511:0] T24;
  wire[7:0] T25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire[29:0] T28;
  wire[27:0] T29;
  wire[25:0] T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire[511:0] T33;
  wire[3:0] T34;
  wire[3:0] T35;
  wire[25:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire T39;
  wire empty;
  wire T40;
  reg  maybe_full;
  wire T41;
  wire T42;
  wire T43;
  wire ptr_match;
  wire T44;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {18{$random}};
    enq_ptr = {1{$random}};
    deq_ptr = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_r_type = T0;
  assign T0 = T1[2'h2:1'h0];
  assign T1 = {T28, T2};
  assign T2 = {T25, T3};
  assign T3 = {T24, T4};
  assign T4 = T5[2'h2:1'h0];
  assign T5 = ram[deq_ptr];
  always @(posedge clk)
    if (do_enq)
      ram[enq_ptr] <= T7;
  assign T7 = T8;
  assign T8 = {T12, T9};
  assign T9 = {T11, T10};
  assign T10 = {io_enq_bits_payload_data, io_enq_bits_payload_r_type};
  assign T11 = {io_enq_bits_payload_client_xact_id, io_enq_bits_payload_master_xact_id};
  assign T12 = {io_enq_bits_header_src, T13};
  assign T13 = {io_enq_bits_header_dst, io_enq_bits_payload_addr};
  assign do_enq = T15 & T14;
  assign T14 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T15 = io_enq_ready & io_enq_valid;
  assign T16 = reset ? 1'h0 : T17;
  assign T17 = do_enq ? T18 : enq_ptr;
  assign T18 = enq_ptr + 1'h1;
  assign T19 = reset ? 1'h0 : T20;
  assign T20 = do_deq ? T21 : deq_ptr;
  assign T21 = deq_ptr + 1'h1;
  assign do_deq = T23 & T22;
  assign T22 = do_flow ^ 1'h1;
  assign T23 = io_deq_ready & io_deq_valid;
  assign T24 = T5[10'h202:2'h3];
  assign T25 = {T27, T26};
  assign T26 = T5[10'h206:10'h203];
  assign T27 = T5[10'h20a:10'h207];
  assign T28 = {T32, T29};
  assign T29 = {T31, T30};
  assign T30 = T5[10'h224:10'h20b];
  assign T31 = T5[10'h226:10'h225];
  assign T32 = T5[10'h228:10'h227];
  assign io_deq_bits_payload_data = T33;
  assign T33 = T1[10'h202:2'h3];
  assign io_deq_bits_payload_master_xact_id = T34;
  assign T34 = T1[10'h206:10'h203];
  assign io_deq_bits_payload_client_xact_id = T35;
  assign T35 = T1[10'h20a:10'h207];
  assign io_deq_bits_payload_addr = T36;
  assign T36 = T1[10'h224:10'h20b];
  assign io_deq_bits_header_dst = T37;
  assign T37 = T1[10'h226:10'h225];
  assign io_deq_bits_header_src = T38;
  assign T38 = T1[10'h228:10'h227];
  assign io_deq_valid = T39;
  assign T39 = empty ^ 1'h1;
  assign empty = ptr_match & T40;
  assign T40 = maybe_full ^ 1'h1;
  assign T41 = reset ? 1'h0 : T42;
  assign T42 = T43 ? do_enq : maybe_full;
  assign T43 = do_enq != do_deq;
  assign ptr_match = enq_ptr == deq_ptr;
  assign io_enq_ready = T44;
  assign T44 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      enq_ptr <= 1'h0;
    end else if(do_enq) begin
      enq_ptr <= T18;
    end
    if(reset) begin
      deq_ptr <= 1'h0;
    end else if(do_deq) begin
      deq_ptr <= T21;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T43) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_10(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [3:0] io_enq_bits_payload_master_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[3:0] io_deq_bits_payload_master_xact_id
);

  wire[3:0] T0;
  wire[7:0] T1;
  wire[5:0] T2;
  wire[3:0] T3;
  wire[7:0] T4;
  reg [7:0] ram [1:0];
  wire[7:0] T5;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[5:0] T8;
  wire do_enq;
  wire T9;
  wire do_flow;
  wire T10;
  reg  enq_ptr;
  wire T11;
  wire T12;
  wire T13;
  reg  deq_ptr;
  wire T14;
  wire T15;
  wire T16;
  wire do_deq;
  wire T17;
  wire T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire[1:0] T22;
  wire T23;
  wire empty;
  wire T24;
  reg  maybe_full;
  wire T25;
  wire T26;
  wire T27;
  wire ptr_match;
  wire T28;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    enq_ptr = {1{$random}};
    deq_ptr = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_master_xact_id = T0;
  assign T0 = T1[2'h3:1'h0];
  assign T1 = {T20, T2};
  assign T2 = {T19, T3};
  assign T3 = T4[2'h3:1'h0];
  assign T4 = ram[deq_ptr];
  always @(posedge clk)
    if (do_enq)
      ram[enq_ptr] <= T6;
  assign T6 = T7;
  assign T7 = {io_enq_bits_header_src, T8};
  assign T8 = {io_enq_bits_header_dst, io_enq_bits_payload_master_xact_id};
  assign do_enq = T10 & T9;
  assign T9 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T10 = io_enq_ready & io_enq_valid;
  assign T11 = reset ? 1'h0 : T12;
  assign T12 = do_enq ? T13 : enq_ptr;
  assign T13 = enq_ptr + 1'h1;
  assign T14 = reset ? 1'h0 : T15;
  assign T15 = do_deq ? T16 : deq_ptr;
  assign T16 = deq_ptr + 1'h1;
  assign do_deq = T18 & T17;
  assign T17 = do_flow ^ 1'h1;
  assign T18 = io_deq_ready & io_deq_valid;
  assign T19 = T4[3'h5:3'h4];
  assign T20 = T4[3'h7:3'h6];
  assign io_deq_bits_header_dst = T21;
  assign T21 = T1[3'h5:3'h4];
  assign io_deq_bits_header_src = T22;
  assign T22 = T1[3'h7:3'h6];
  assign io_deq_valid = T23;
  assign T23 = empty ^ 1'h1;
  assign empty = ptr_match & T24;
  assign T24 = maybe_full ^ 1'h1;
  assign T25 = reset ? 1'h0 : T26;
  assign T26 = T27 ? do_enq : maybe_full;
  assign T27 = do_enq != do_deq;
  assign ptr_match = enq_ptr == deq_ptr;
  assign io_enq_ready = T28;
  assign T28 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      enq_ptr <= 1'h0;
    end else if(do_enq) begin
      enq_ptr <= T13;
    end
    if(reset) begin
      deq_ptr <= 1'h0;
    end else if(do_deq) begin
      deq_ptr <= T16;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T27) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_11(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [511:0] io_enq_bits_payload_data,
    input [3:0] io_enq_bits_payload_client_xact_id,
    input [3:0] io_enq_bits_payload_master_xact_id,
    input [3:0] io_enq_bits_payload_g_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[511:0] io_deq_bits_payload_data,
    output[3:0] io_deq_bits_payload_client_xact_id,
    output[3:0] io_deq_bits_payload_master_xact_id,
    output[3:0] io_deq_bits_payload_g_type
);

  wire[3:0] T0;
  wire[527:0] T1;
  wire[11:0] T2;
  wire[7:0] T3;
  wire[3:0] T4;
  wire[527:0] T5;
  reg [527:0] ram [0:0];
  wire[527:0] T6;
  wire[527:0] T7;
  wire[527:0] T8;
  wire[11:0] T9;
  wire[7:0] T10;
  wire[515:0] T11;
  wire[513:0] T12;
  wire do_enq;
  wire T13;
  wire do_flow;
  wire T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[515:0] T17;
  wire[513:0] T18;
  wire[511:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire[3:0] T22;
  wire[3:0] T23;
  wire[511:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire T27;
  wire empty;
  reg  maybe_full;
  wire T28;
  wire T29;
  wire T30;
  wire do_deq;
  wire T31;
  wire T32;
  wire T33;
  wire T34;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {17{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_g_type = T0;
  assign T0 = T1[2'h3:1'h0];
  assign T1 = {T17, T2};
  assign T2 = {T16, T3};
  assign T3 = {T15, T4};
  assign T4 = T5[2'h3:1'h0];
  assign T5 = ram[1'h0];
  always @(posedge clk)
    if (do_enq)
      ram[1'h0] <= T7;
  assign T7 = T8;
  assign T8 = {T11, T9};
  assign T9 = {io_enq_bits_payload_client_xact_id, T10};
  assign T10 = {io_enq_bits_payload_master_xact_id, io_enq_bits_payload_g_type};
  assign T11 = {io_enq_bits_header_src, T12};
  assign T12 = {io_enq_bits_header_dst, io_enq_bits_payload_data};
  assign do_enq = T14 & T13;
  assign T13 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T14 = io_enq_ready & io_enq_valid;
  assign T15 = T5[3'h7:3'h4];
  assign T16 = T5[4'hb:4'h8];
  assign T17 = {T21, T18};
  assign T18 = {T20, T19};
  assign T19 = T5[10'h20b:4'hc];
  assign T20 = T5[10'h20d:10'h20c];
  assign T21 = T5[10'h20f:10'h20e];
  assign io_deq_bits_payload_master_xact_id = T22;
  assign T22 = T1[3'h7:3'h4];
  assign io_deq_bits_payload_client_xact_id = T23;
  assign T23 = T1[4'hb:4'h8];
  assign io_deq_bits_payload_data = T24;
  assign T24 = T1[10'h20b:4'hc];
  assign io_deq_bits_header_dst = T25;
  assign T25 = T1[10'h20d:10'h20c];
  assign io_deq_bits_header_src = T26;
  assign T26 = T1[10'h20f:10'h20e];
  assign io_deq_valid = T27;
  assign T27 = empty ^ 1'h1;
  assign empty = maybe_full ^ 1'h1;
  assign T28 = reset ? 1'h0 : T29;
  assign T29 = T30 ? do_enq : maybe_full;
  assign T30 = do_enq != do_deq;
  assign do_deq = T32 & T31;
  assign T31 = do_flow ^ 1'h1;
  assign T32 = io_deq_ready & io_deq_valid;
  assign io_enq_ready = T33;
  assign T33 = T34 | io_deq_ready;
  assign T34 = maybe_full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T30) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_12(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [3:0] io_enq_bits_payload_master_xact_id,
    input [1:0] io_enq_bits_payload_p_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[3:0] io_deq_bits_payload_master_xact_id,
    output[1:0] io_deq_bits_payload_p_type
);

  wire[1:0] T0;
  wire[35:0] T1;
  wire[31:0] T2;
  wire[5:0] T3;
  wire[1:0] T4;
  wire[35:0] T5;
  reg [35:0] ram [1:0];
  wire[35:0] T6;
  wire[35:0] T7;
  wire[35:0] T8;
  wire[31:0] T9;
  wire[5:0] T10;
  wire[3:0] T11;
  wire do_enq;
  wire T12;
  wire do_flow;
  wire T13;
  reg  enq_ptr;
  wire T14;
  wire T15;
  wire T16;
  reg  deq_ptr;
  wire T17;
  wire T18;
  wire T19;
  wire do_deq;
  wire T20;
  wire T21;
  wire[3:0] T22;
  wire[25:0] T23;
  wire[3:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire[3:0] T27;
  wire[25:0] T28;
  wire[1:0] T29;
  wire[1:0] T30;
  wire T31;
  wire empty;
  wire T32;
  reg  maybe_full;
  wire T33;
  wire T34;
  wire T35;
  wire ptr_match;
  wire T36;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
    enq_ptr = {1{$random}};
    deq_ptr = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_p_type = T0;
  assign T0 = T1[1'h1:1'h0];
  assign T1 = {T24, T2};
  assign T2 = {T23, T3};
  assign T3 = {T22, T4};
  assign T4 = T5[1'h1:1'h0];
  assign T5 = ram[deq_ptr];
  always @(posedge clk)
    if (do_enq)
      ram[enq_ptr] <= T7;
  assign T7 = T8;
  assign T8 = {T11, T9};
  assign T9 = {io_enq_bits_payload_addr, T10};
  assign T10 = {io_enq_bits_payload_master_xact_id, io_enq_bits_payload_p_type};
  assign T11 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign do_enq = T13 & T12;
  assign T12 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T13 = io_enq_ready & io_enq_valid;
  assign T14 = reset ? 1'h0 : T15;
  assign T15 = do_enq ? T16 : enq_ptr;
  assign T16 = enq_ptr + 1'h1;
  assign T17 = reset ? 1'h0 : T18;
  assign T18 = do_deq ? T19 : deq_ptr;
  assign T19 = deq_ptr + 1'h1;
  assign do_deq = T21 & T20;
  assign T20 = do_flow ^ 1'h1;
  assign T21 = io_deq_ready & io_deq_valid;
  assign T22 = T5[3'h5:2'h2];
  assign T23 = T5[5'h1f:3'h6];
  assign T24 = {T26, T25};
  assign T25 = T5[6'h21:6'h20];
  assign T26 = T5[6'h23:6'h22];
  assign io_deq_bits_payload_master_xact_id = T27;
  assign T27 = T1[3'h5:2'h2];
  assign io_deq_bits_payload_addr = T28;
  assign T28 = T1[5'h1f:3'h6];
  assign io_deq_bits_header_dst = T29;
  assign T29 = T1[6'h21:6'h20];
  assign io_deq_bits_header_src = T30;
  assign T30 = T1[6'h23:6'h22];
  assign io_deq_valid = T31;
  assign T31 = empty ^ 1'h1;
  assign empty = ptr_match & T32;
  assign T32 = maybe_full ^ 1'h1;
  assign T33 = reset ? 1'h0 : T34;
  assign T34 = T35 ? do_enq : maybe_full;
  assign T35 = do_enq != do_deq;
  assign ptr_match = enq_ptr == deq_ptr;
  assign io_enq_ready = T36;
  assign T36 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      enq_ptr <= 1'h0;
    end else if(do_enq) begin
      enq_ptr <= T16;
    end
    if(reset) begin
      deq_ptr <= 1'h0;
    end else if(do_deq) begin
      deq_ptr <= T19;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T35) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module FPGAUncore(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    //output io_host_debug_stats_pcr
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    output io_mem_resp_ready,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag,
    output io_tiles_0_acquire_ready,
    input  io_tiles_0_acquire_valid,
    input [1:0] io_tiles_0_acquire_bits_header_src,
    input [1:0] io_tiles_0_acquire_bits_header_dst,
    input [25:0] io_tiles_0_acquire_bits_payload_addr,
    input [3:0] io_tiles_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_tiles_0_acquire_bits_payload_data,
    input [2:0] io_tiles_0_acquire_bits_payload_a_type,
    input [5:0] io_tiles_0_acquire_bits_payload_write_mask,
    input [2:0] io_tiles_0_acquire_bits_payload_subword_addr,
    input [3:0] io_tiles_0_acquire_bits_payload_atomic_opcode,
    input  io_tiles_0_grant_ready,
    output io_tiles_0_grant_valid,
    output[1:0] io_tiles_0_grant_bits_header_src,
    output[1:0] io_tiles_0_grant_bits_header_dst,
    output[511:0] io_tiles_0_grant_bits_payload_data,
    output[3:0] io_tiles_0_grant_bits_payload_client_xact_id,
    output[3:0] io_tiles_0_grant_bits_payload_master_xact_id,
    output[3:0] io_tiles_0_grant_bits_payload_g_type,
    output io_tiles_0_finish_ready,
    input  io_tiles_0_finish_valid,
    input [1:0] io_tiles_0_finish_bits_header_src,
    input [1:0] io_tiles_0_finish_bits_header_dst,
    input [3:0] io_tiles_0_finish_bits_payload_master_xact_id,
    input  io_tiles_0_probe_ready,
    output io_tiles_0_probe_valid,
    output[1:0] io_tiles_0_probe_bits_header_src,
    output[1:0] io_tiles_0_probe_bits_header_dst,
    output[25:0] io_tiles_0_probe_bits_payload_addr,
    output[3:0] io_tiles_0_probe_bits_payload_master_xact_id,
    output[1:0] io_tiles_0_probe_bits_payload_p_type,
    output io_tiles_0_release_ready,
    input  io_tiles_0_release_valid,
    input [1:0] io_tiles_0_release_bits_header_src,
    input [1:0] io_tiles_0_release_bits_header_dst,
    input [25:0] io_tiles_0_release_bits_payload_addr,
    input [3:0] io_tiles_0_release_bits_payload_client_xact_id,
    input [3:0] io_tiles_0_release_bits_payload_master_xact_id,
    input [511:0] io_tiles_0_release_bits_payload_data,
    input [2:0] io_tiles_0_release_bits_payload_r_type,
    output io_htif_0_reset,
    //output io_htif_0_id
    input  io_htif_0_pcr_req_ready,
    output io_htif_0_pcr_req_valid,
    output io_htif_0_pcr_req_bits_rw,
    output[4:0] io_htif_0_pcr_req_bits_addr,
    output[63:0] io_htif_0_pcr_req_bits_data,
    output io_htif_0_pcr_rep_ready,
    input  io_htif_0_pcr_rep_valid,
    input [63:0] io_htif_0_pcr_rep_bits,
    output io_htif_0_ipi_req_ready,
    input  io_htif_0_ipi_req_valid,
    input  io_htif_0_ipi_req_bits,
    input  io_htif_0_ipi_rep_ready,
    output io_htif_0_ipi_rep_valid,
    output io_htif_0_ipi_rep_bits,
    input  io_htif_0_debug_stats_pcr,
    input  io_incoherent_0
);

  wire htif_io_mem_probe_ready;
  wire[1:0] outmemsys_io_htif_probe_bits_payload_p_type;
  wire[3:0] outmemsys_io_htif_probe_bits_payload_master_xact_id;
  wire[25:0] outmemsys_io_htif_probe_bits_payload_addr;
  wire[1:0] outmemsys_io_htif_probe_bits_header_dst;
  wire[1:0] outmemsys_io_htif_probe_bits_header_src;
  wire outmemsys_io_htif_probe_valid;
  wire htif_io_mem_grant_ready;
  wire[3:0] outmemsys_io_htif_grant_bits_payload_g_type;
  wire[3:0] outmemsys_io_htif_grant_bits_payload_master_xact_id;
  wire[3:0] outmemsys_io_htif_grant_bits_payload_client_xact_id;
  wire[511:0] outmemsys_io_htif_grant_bits_payload_data;
  wire[1:0] outmemsys_io_htif_grant_bits_header_dst;
  wire[1:0] outmemsys_io_htif_grant_bits_header_src;
  wire outmemsys_io_htif_grant_valid;
  wire outmemsys_io_htif_finish_ready;
  wire[3:0] T0;
  wire[3:0] htif_io_mem_finish_bits_payload_master_xact_id;
  wire[1:0] T1;
  wire[1:0] htif_io_mem_finish_bits_header_dst;
  wire[1:0] T2;
  wire T3;
  wire htif_io_mem_finish_valid;
  wire outmemsys_io_htif_release_ready;
  wire[2:0] T4;
  wire[2:0] htif_io_mem_release_bits_payload_r_type;
  wire[511:0] T5;
  wire[511:0] htif_io_mem_release_bits_payload_data;
  wire[3:0] T6;
  wire[3:0] htif_io_mem_release_bits_payload_master_xact_id;
  wire[3:0] T7;
  wire[3:0] htif_io_mem_release_bits_payload_client_xact_id;
  wire[25:0] T8;
  wire[25:0] htif_io_mem_release_bits_payload_addr;
  wire[1:0] T9;
  wire[1:0] T10;
  wire T11;
  wire htif_io_mem_release_valid;
  wire outmemsys_io_htif_acquire_ready;
  wire[3:0] T12;
  wire[3:0] htif_io_mem_acquire_bits_payload_atomic_opcode;
  wire[2:0] T13;
  wire[2:0] htif_io_mem_acquire_bits_payload_subword_addr;
  wire[5:0] T14;
  wire[5:0] htif_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] T15;
  wire[2:0] htif_io_mem_acquire_bits_payload_a_type;
  wire[511:0] T16;
  wire[511:0] htif_io_mem_acquire_bits_payload_data;
  wire[3:0] T17;
  wire[3:0] htif_io_mem_acquire_bits_payload_client_xact_id;
  wire[25:0] T18;
  wire[25:0] htif_io_mem_acquire_bits_payload_addr;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire htif_io_mem_acquire_valid;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_payload_p_type;
  wire[3:0] outmemsys_io_tiles_0_probe_bits_payload_master_xact_id;
  wire[25:0] outmemsys_io_tiles_0_probe_bits_payload_addr;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_header_dst;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_header_src;
  wire outmemsys_io_tiles_0_probe_valid;
  wire[3:0] outmemsys_io_tiles_0_grant_bits_payload_g_type;
  wire[3:0] outmemsys_io_tiles_0_grant_bits_payload_master_xact_id;
  wire[3:0] outmemsys_io_tiles_0_grant_bits_payload_client_xact_id;
  wire[511:0] outmemsys_io_tiles_0_grant_bits_payload_data;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_header_dst;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_header_src;
  wire outmemsys_io_tiles_0_grant_valid;
  wire outmemsys_io_tiles_0_finish_ready;
  wire[3:0] T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire outmemsys_io_tiles_0_release_ready;
  wire[2:0] T26;
  wire[511:0] T27;
  wire[3:0] T28;
  wire[3:0] T29;
  wire[25:0] T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire outmemsys_io_tiles_0_acquire_ready;
  wire[3:0] T34;
  wire[2:0] T35;
  wire[5:0] T36;
  wire[2:0] T37;
  wire[511:0] T38;
  wire[3:0] T39;
  wire[25:0] T40;
  wire[1:0] T41;
  wire[1:0] T42;
  wire T43;
  wire[2:0] Queue_6_io_deq_bits_payload_r_type;
  wire[511:0] Queue_6_io_deq_bits_payload_data;
  wire[3:0] Queue_6_io_deq_bits_payload_master_xact_id;
  wire[3:0] Queue_6_io_deq_bits_payload_client_xact_id;
  wire[25:0] Queue_6_io_deq_bits_payload_addr;
  wire[1:0] Queue_6_io_deq_bits_header_dst;
  wire[1:0] Queue_6_io_deq_bits_header_src;
  wire Queue_6_io_deq_valid;
  wire Queue_9_io_enq_ready;
  wire[3:0] Queue_7_io_deq_bits_payload_master_xact_id;
  wire[1:0] Queue_7_io_deq_bits_header_dst;
  wire[1:0] Queue_7_io_deq_bits_header_src;
  wire Queue_7_io_deq_valid;
  wire Queue_8_io_enq_ready;
  wire[3:0] Queue_5_io_deq_bits_payload_atomic_opcode;
  wire[2:0] Queue_5_io_deq_bits_payload_subword_addr;
  wire[5:0] Queue_5_io_deq_bits_payload_write_mask;
  wire[2:0] Queue_5_io_deq_bits_payload_a_type;
  wire[511:0] Queue_5_io_deq_bits_payload_data;
  wire[3:0] Queue_5_io_deq_bits_payload_client_xact_id;
  wire[25:0] Queue_5_io_deq_bits_payload_addr;
  wire[1:0] Queue_5_io_deq_bits_header_dst;
  wire[1:0] Queue_5_io_deq_bits_header_src;
  wire Queue_5_io_deq_valid;
  wire[2:0] Queue_1_io_deq_bits_payload_r_type;
  wire[511:0] Queue_1_io_deq_bits_payload_data;
  wire[3:0] Queue_1_io_deq_bits_payload_master_xact_id;
  wire[3:0] Queue_1_io_deq_bits_payload_client_xact_id;
  wire[25:0] Queue_1_io_deq_bits_payload_addr;
  wire[1:0] Queue_1_io_deq_bits_header_dst;
  wire[1:0] Queue_1_io_deq_bits_header_src;
  wire Queue_1_io_deq_valid;
  wire Queue_4_io_enq_ready;
  wire[3:0] Queue_2_io_deq_bits_payload_master_xact_id;
  wire[1:0] Queue_2_io_deq_bits_header_dst;
  wire[1:0] Queue_2_io_deq_bits_header_src;
  wire Queue_2_io_deq_valid;
  wire Queue_3_io_enq_ready;
  wire[3:0] Queue_0_io_deq_bits_payload_atomic_opcode;
  wire[2:0] Queue_0_io_deq_bits_payload_subword_addr;
  wire[5:0] Queue_0_io_deq_bits_payload_write_mask;
  wire[2:0] Queue_0_io_deq_bits_payload_a_type;
  wire[511:0] Queue_0_io_deq_bits_payload_data;
  wire[3:0] Queue_0_io_deq_bits_payload_client_xact_id;
  wire[25:0] Queue_0_io_deq_bits_payload_addr;
  wire[1:0] Queue_0_io_deq_bits_header_dst;
  wire[1:0] Queue_0_io_deq_bits_header_src;
  wire Queue_0_io_deq_valid;
  wire T44;
  wire Queue_6_io_enq_ready;
  wire[1:0] Queue_9_io_deq_bits_payload_p_type;
  wire[3:0] Queue_9_io_deq_bits_payload_master_xact_id;
  wire[25:0] Queue_9_io_deq_bits_payload_addr;
  wire[1:0] Queue_9_io_deq_bits_header_dst;
  wire[1:0] Queue_9_io_deq_bits_header_src;
  wire Queue_9_io_deq_valid;
  wire T45;
  wire Queue_7_io_enq_ready;
  wire[3:0] Queue_8_io_deq_bits_payload_g_type;
  wire[3:0] Queue_8_io_deq_bits_payload_master_xact_id;
  wire[3:0] Queue_8_io_deq_bits_payload_client_xact_id;
  wire[511:0] Queue_8_io_deq_bits_payload_data;
  wire[1:0] Queue_8_io_deq_bits_header_dst;
  wire[1:0] Queue_8_io_deq_bits_header_src;
  wire Queue_8_io_deq_valid;
  wire T46;
  wire Queue_5_io_enq_ready;
  wire htif_io_cpu_0_ipi_rep_valid;
  wire htif_io_cpu_0_ipi_req_ready;
  wire htif_io_cpu_0_pcr_rep_ready;
  wire[63:0] htif_io_cpu_0_pcr_req_bits_data;
  wire[4:0] htif_io_cpu_0_pcr_req_bits_addr;
  wire htif_io_cpu_0_pcr_req_bits_rw;
  wire htif_io_cpu_0_pcr_req_valid;
  wire htif_io_cpu_0_reset;
  wire T47;
  wire Queue_1_io_enq_ready;
  wire[1:0] Queue_4_io_deq_bits_payload_p_type;
  wire[3:0] Queue_4_io_deq_bits_payload_master_xact_id;
  wire[25:0] Queue_4_io_deq_bits_payload_addr;
  wire[1:0] Queue_4_io_deq_bits_header_dst;
  wire[1:0] Queue_4_io_deq_bits_header_src;
  wire Queue_4_io_deq_valid;
  wire T48;
  wire Queue_2_io_enq_ready;
  wire[3:0] Queue_3_io_deq_bits_payload_g_type;
  wire[3:0] Queue_3_io_deq_bits_payload_master_xact_id;
  wire[3:0] Queue_3_io_deq_bits_payload_client_xact_id;
  wire[511:0] Queue_3_io_deq_bits_payload_data;
  wire[1:0] Queue_3_io_deq_bits_header_dst;
  wire[1:0] Queue_3_io_deq_bits_header_src;
  wire Queue_3_io_deq_valid;
  wire T49;
  wire Queue_0_io_enq_ready;
  wire outmemsys_io_mem_resp_ready;
  wire[127:0] outmemsys_io_mem_req_data_bits_data;
  wire outmemsys_io_mem_req_data_valid;
  wire outmemsys_io_mem_req_cmd_bits_rw;
  wire[4:0] outmemsys_io_mem_req_cmd_bits_tag;
  wire[25:0] outmemsys_io_mem_req_cmd_bits_addr;
  wire outmemsys_io_mem_req_cmd_valid;
  wire[15:0] htif_io_host_out_bits;
  wire htif_io_host_out_valid;
  wire htif_io_host_in_ready;


  assign T0 = htif_io_mem_finish_bits_payload_master_xact_id;
  assign T1 = htif_io_mem_finish_bits_header_dst;
  assign T2 = 2'h1;
  assign T3 = htif_io_mem_finish_valid;
  assign T4 = htif_io_mem_release_bits_payload_r_type;
  assign T5 = htif_io_mem_release_bits_payload_data;
  assign T6 = htif_io_mem_release_bits_payload_master_xact_id;
  assign T7 = htif_io_mem_release_bits_payload_client_xact_id;
  assign T8 = htif_io_mem_release_bits_payload_addr;
  assign T9 = 2'h0;
  assign T10 = 2'h1;
  assign T11 = htif_io_mem_release_valid;
  assign T12 = htif_io_mem_acquire_bits_payload_atomic_opcode;
  assign T13 = htif_io_mem_acquire_bits_payload_subword_addr;
  assign T14 = htif_io_mem_acquire_bits_payload_write_mask;
  assign T15 = htif_io_mem_acquire_bits_payload_a_type;
  assign T16 = htif_io_mem_acquire_bits_payload_data;
  assign T17 = htif_io_mem_acquire_bits_payload_client_xact_id;
  assign T18 = htif_io_mem_acquire_bits_payload_addr;
  assign T19 = 2'h0;
  assign T20 = 2'h1;
  assign T21 = htif_io_mem_acquire_valid;
  assign T22 = io_tiles_0_finish_bits_payload_master_xact_id;
  assign T23 = io_tiles_0_finish_bits_header_dst;
  assign T24 = 2'h0;
  assign T25 = io_tiles_0_finish_valid;
  assign T26 = io_tiles_0_release_bits_payload_r_type;
  assign T27 = io_tiles_0_release_bits_payload_data;
  assign T28 = io_tiles_0_release_bits_payload_master_xact_id;
  assign T29 = io_tiles_0_release_bits_payload_client_xact_id;
  assign T30 = io_tiles_0_release_bits_payload_addr;
  assign T31 = 2'h0;
  assign T32 = 2'h0;
  assign T33 = io_tiles_0_release_valid;
  assign T34 = io_tiles_0_acquire_bits_payload_atomic_opcode;
  assign T35 = io_tiles_0_acquire_bits_payload_subword_addr;
  assign T36 = io_tiles_0_acquire_bits_payload_write_mask;
  assign T37 = io_tiles_0_acquire_bits_payload_a_type;
  assign T38 = io_tiles_0_acquire_bits_payload_data;
  assign T39 = io_tiles_0_acquire_bits_payload_client_xact_id;
  assign T40 = io_tiles_0_acquire_bits_payload_addr;
  assign T41 = 2'h0;
  assign T42 = 2'h0;
  assign T43 = io_tiles_0_acquire_valid;
  assign T44 = Queue_6_io_enq_ready;
  assign T45 = Queue_7_io_enq_ready;
  assign T46 = Queue_5_io_enq_ready;
  assign io_htif_0_ipi_rep_valid = htif_io_cpu_0_ipi_rep_valid;
  assign io_htif_0_ipi_req_ready = htif_io_cpu_0_ipi_req_ready;
  assign io_htif_0_pcr_rep_ready = htif_io_cpu_0_pcr_rep_ready;
  assign io_htif_0_pcr_req_bits_data = htif_io_cpu_0_pcr_req_bits_data;
  assign io_htif_0_pcr_req_bits_addr = htif_io_cpu_0_pcr_req_bits_addr;
  assign io_htif_0_pcr_req_bits_rw = htif_io_cpu_0_pcr_req_bits_rw;
  assign io_htif_0_pcr_req_valid = htif_io_cpu_0_pcr_req_valid;
  assign io_htif_0_reset = htif_io_cpu_0_reset;
  assign io_tiles_0_release_ready = T47;
  assign T47 = Queue_1_io_enq_ready;
  assign io_tiles_0_probe_bits_payload_p_type = Queue_4_io_deq_bits_payload_p_type;
  assign io_tiles_0_probe_bits_payload_master_xact_id = Queue_4_io_deq_bits_payload_master_xact_id;
  assign io_tiles_0_probe_bits_payload_addr = Queue_4_io_deq_bits_payload_addr;
  assign io_tiles_0_probe_bits_header_dst = Queue_4_io_deq_bits_header_dst;
  assign io_tiles_0_probe_bits_header_src = Queue_4_io_deq_bits_header_src;
  assign io_tiles_0_probe_valid = Queue_4_io_deq_valid;
  assign io_tiles_0_finish_ready = T48;
  assign T48 = Queue_2_io_enq_ready;
  assign io_tiles_0_grant_bits_payload_g_type = Queue_3_io_deq_bits_payload_g_type;
  assign io_tiles_0_grant_bits_payload_master_xact_id = Queue_3_io_deq_bits_payload_master_xact_id;
  assign io_tiles_0_grant_bits_payload_client_xact_id = Queue_3_io_deq_bits_payload_client_xact_id;
  assign io_tiles_0_grant_bits_payload_data = Queue_3_io_deq_bits_payload_data;
  assign io_tiles_0_grant_bits_header_dst = Queue_3_io_deq_bits_header_dst;
  assign io_tiles_0_grant_bits_header_src = Queue_3_io_deq_bits_header_src;
  assign io_tiles_0_grant_valid = Queue_3_io_deq_valid;
  assign io_tiles_0_acquire_ready = T49;
  assign T49 = Queue_0_io_enq_ready;
  assign io_mem_resp_ready = outmemsys_io_mem_resp_ready;
  assign io_mem_req_data_bits_data = outmemsys_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = outmemsys_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = outmemsys_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = outmemsys_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = outmemsys_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = outmemsys_io_mem_req_cmd_valid;
  assign io_host_out_bits = htif_io_host_out_bits;
  assign io_host_out_valid = htif_io_host_out_valid;
  assign io_host_in_ready = htif_io_host_in_ready;
  HTIF htif(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( htif_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( htif_io_host_out_valid ),
       .io_host_out_bits( htif_io_host_out_bits ),
       //.io_host_debug_stats_pcr(  )
       .io_cpu_0_reset( htif_io_cpu_0_reset ),
       //.io_cpu_0_id(  )
       .io_cpu_0_pcr_req_ready( io_htif_0_pcr_req_ready ),
       .io_cpu_0_pcr_req_valid( htif_io_cpu_0_pcr_req_valid ),
       .io_cpu_0_pcr_req_bits_rw( htif_io_cpu_0_pcr_req_bits_rw ),
       .io_cpu_0_pcr_req_bits_addr( htif_io_cpu_0_pcr_req_bits_addr ),
       .io_cpu_0_pcr_req_bits_data( htif_io_cpu_0_pcr_req_bits_data ),
       .io_cpu_0_pcr_rep_ready( htif_io_cpu_0_pcr_rep_ready ),
       .io_cpu_0_pcr_rep_valid( io_htif_0_pcr_rep_valid ),
       .io_cpu_0_pcr_rep_bits( io_htif_0_pcr_rep_bits ),
       .io_cpu_0_ipi_req_ready( htif_io_cpu_0_ipi_req_ready ),
       .io_cpu_0_ipi_req_valid( io_htif_0_ipi_req_valid ),
       .io_cpu_0_ipi_req_bits( io_htif_0_ipi_req_bits ),
       .io_cpu_0_ipi_rep_ready( io_htif_0_ipi_rep_ready ),
       .io_cpu_0_ipi_rep_valid( htif_io_cpu_0_ipi_rep_valid ),
       //.io_cpu_0_ipi_rep_bits(  )
       .io_cpu_0_debug_stats_pcr( io_htif_0_debug_stats_pcr ),
       .io_mem_acquire_ready( T46 ),
       .io_mem_acquire_valid( htif_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( htif_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( htif_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( htif_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( htif_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( htif_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( htif_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( htif_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( htif_io_mem_grant_ready ),
       .io_mem_grant_valid( Queue_8_io_deq_valid ),
       .io_mem_grant_bits_header_src( Queue_8_io_deq_bits_header_src ),
       .io_mem_grant_bits_header_dst( Queue_8_io_deq_bits_header_dst ),
       .io_mem_grant_bits_payload_data( Queue_8_io_deq_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( Queue_8_io_deq_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( Queue_8_io_deq_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( Queue_8_io_deq_bits_payload_g_type ),
       .io_mem_finish_ready( T45 ),
       .io_mem_finish_valid( htif_io_mem_finish_valid ),
       //.io_mem_finish_bits_header_src(  )
       .io_mem_finish_bits_header_dst( htif_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( htif_io_mem_finish_bits_payload_master_xact_id ),
       .io_mem_probe_ready( htif_io_mem_probe_ready ),
       .io_mem_probe_valid( Queue_9_io_deq_valid ),
       .io_mem_probe_bits_header_src( Queue_9_io_deq_bits_header_src ),
       .io_mem_probe_bits_header_dst( Queue_9_io_deq_bits_header_dst ),
       .io_mem_probe_bits_payload_addr( Queue_9_io_deq_bits_payload_addr ),
       .io_mem_probe_bits_payload_master_xact_id( Queue_9_io_deq_bits_payload_master_xact_id ),
       .io_mem_probe_bits_payload_p_type( Queue_9_io_deq_bits_payload_p_type ),
       .io_mem_release_ready( T44 ),
       .io_mem_release_valid( htif_io_mem_release_valid ),
       //.io_mem_release_bits_header_src(  )
       //.io_mem_release_bits_header_dst(  )
       .io_mem_release_bits_payload_addr( htif_io_mem_release_bits_payload_addr ),
       .io_mem_release_bits_payload_client_xact_id( htif_io_mem_release_bits_payload_client_xact_id ),
       .io_mem_release_bits_payload_master_xact_id( htif_io_mem_release_bits_payload_master_xact_id ),
       .io_mem_release_bits_payload_data( htif_io_mem_release_bits_payload_data ),
       .io_mem_release_bits_payload_r_type( htif_io_mem_release_bits_payload_r_type )
       //.io_scr_rdata_63(  )
       //.io_scr_rdata_62(  )
       //.io_scr_rdata_61(  )
       //.io_scr_rdata_60(  )
       //.io_scr_rdata_59(  )
       //.io_scr_rdata_58(  )
       //.io_scr_rdata_57(  )
       //.io_scr_rdata_56(  )
       //.io_scr_rdata_55(  )
       //.io_scr_rdata_54(  )
       //.io_scr_rdata_53(  )
       //.io_scr_rdata_52(  )
       //.io_scr_rdata_51(  )
       //.io_scr_rdata_50(  )
       //.io_scr_rdata_49(  )
       //.io_scr_rdata_48(  )
       //.io_scr_rdata_47(  )
       //.io_scr_rdata_46(  )
       //.io_scr_rdata_45(  )
       //.io_scr_rdata_44(  )
       //.io_scr_rdata_43(  )
       //.io_scr_rdata_42(  )
       //.io_scr_rdata_41(  )
       //.io_scr_rdata_40(  )
       //.io_scr_rdata_39(  )
       //.io_scr_rdata_38(  )
       //.io_scr_rdata_37(  )
       //.io_scr_rdata_36(  )
       //.io_scr_rdata_35(  )
       //.io_scr_rdata_34(  )
       //.io_scr_rdata_33(  )
       //.io_scr_rdata_32(  )
       //.io_scr_rdata_31(  )
       //.io_scr_rdata_30(  )
       //.io_scr_rdata_29(  )
       //.io_scr_rdata_28(  )
       //.io_scr_rdata_27(  )
       //.io_scr_rdata_26(  )
       //.io_scr_rdata_25(  )
       //.io_scr_rdata_24(  )
       //.io_scr_rdata_23(  )
       //.io_scr_rdata_22(  )
       //.io_scr_rdata_21(  )
       //.io_scr_rdata_20(  )
       //.io_scr_rdata_19(  )
       //.io_scr_rdata_18(  )
       //.io_scr_rdata_17(  )
       //.io_scr_rdata_16(  )
       //.io_scr_rdata_15(  )
       //.io_scr_rdata_14(  )
       //.io_scr_rdata_13(  )
       //.io_scr_rdata_12(  )
       //.io_scr_rdata_11(  )
       //.io_scr_rdata_10(  )
       //.io_scr_rdata_9(  )
       //.io_scr_rdata_8(  )
       //.io_scr_rdata_7(  )
       //.io_scr_rdata_6(  )
       //.io_scr_rdata_5(  )
       //.io_scr_rdata_4(  )
       //.io_scr_rdata_3(  )
       //.io_scr_rdata_2(  )
       //.io_scr_rdata_1(  )
       //.io_scr_rdata_0(  )
       //.io_scr_wen(  )
       //.io_scr_waddr(  )
       //.io_scr_wdata(  )
  );
  `ifndef SYNTHESIS
    assign htif.io_mem_release_bits_payload_addr = {1{$random}};
    assign htif.io_mem_release_bits_payload_client_xact_id = {1{$random}};
    assign htif.io_mem_release_bits_payload_master_xact_id = {1{$random}};
    assign htif.io_mem_release_bits_payload_data = {16{$random}};
    assign htif.io_mem_release_bits_payload_r_type = {1{$random}};
    assign htif.io_scr_rdata_63 = {2{$random}};
    assign htif.io_scr_rdata_62 = {2{$random}};
    assign htif.io_scr_rdata_61 = {2{$random}};
    assign htif.io_scr_rdata_60 = {2{$random}};
    assign htif.io_scr_rdata_59 = {2{$random}};
    assign htif.io_scr_rdata_58 = {2{$random}};
    assign htif.io_scr_rdata_57 = {2{$random}};
    assign htif.io_scr_rdata_56 = {2{$random}};
    assign htif.io_scr_rdata_55 = {2{$random}};
    assign htif.io_scr_rdata_54 = {2{$random}};
    assign htif.io_scr_rdata_53 = {2{$random}};
    assign htif.io_scr_rdata_52 = {2{$random}};
    assign htif.io_scr_rdata_51 = {2{$random}};
    assign htif.io_scr_rdata_50 = {2{$random}};
    assign htif.io_scr_rdata_49 = {2{$random}};
    assign htif.io_scr_rdata_48 = {2{$random}};
    assign htif.io_scr_rdata_47 = {2{$random}};
    assign htif.io_scr_rdata_46 = {2{$random}};
    assign htif.io_scr_rdata_45 = {2{$random}};
    assign htif.io_scr_rdata_44 = {2{$random}};
    assign htif.io_scr_rdata_43 = {2{$random}};
    assign htif.io_scr_rdata_42 = {2{$random}};
    assign htif.io_scr_rdata_41 = {2{$random}};
    assign htif.io_scr_rdata_40 = {2{$random}};
    assign htif.io_scr_rdata_39 = {2{$random}};
    assign htif.io_scr_rdata_38 = {2{$random}};
    assign htif.io_scr_rdata_37 = {2{$random}};
    assign htif.io_scr_rdata_36 = {2{$random}};
    assign htif.io_scr_rdata_35 = {2{$random}};
    assign htif.io_scr_rdata_34 = {2{$random}};
    assign htif.io_scr_rdata_33 = {2{$random}};
    assign htif.io_scr_rdata_32 = {2{$random}};
    assign htif.io_scr_rdata_31 = {2{$random}};
    assign htif.io_scr_rdata_30 = {2{$random}};
    assign htif.io_scr_rdata_29 = {2{$random}};
    assign htif.io_scr_rdata_28 = {2{$random}};
    assign htif.io_scr_rdata_27 = {2{$random}};
    assign htif.io_scr_rdata_26 = {2{$random}};
    assign htif.io_scr_rdata_25 = {2{$random}};
    assign htif.io_scr_rdata_24 = {2{$random}};
    assign htif.io_scr_rdata_23 = {2{$random}};
    assign htif.io_scr_rdata_22 = {2{$random}};
    assign htif.io_scr_rdata_21 = {2{$random}};
    assign htif.io_scr_rdata_20 = {2{$random}};
    assign htif.io_scr_rdata_19 = {2{$random}};
    assign htif.io_scr_rdata_18 = {2{$random}};
    assign htif.io_scr_rdata_17 = {2{$random}};
    assign htif.io_scr_rdata_16 = {2{$random}};
    assign htif.io_scr_rdata_15 = {2{$random}};
    assign htif.io_scr_rdata_14 = {2{$random}};
    assign htif.io_scr_rdata_13 = {2{$random}};
    assign htif.io_scr_rdata_12 = {2{$random}};
    assign htif.io_scr_rdata_11 = {2{$random}};
    assign htif.io_scr_rdata_10 = {2{$random}};
    assign htif.io_scr_rdata_9 = {2{$random}};
    assign htif.io_scr_rdata_8 = {2{$random}};
    assign htif.io_scr_rdata_7 = {2{$random}};
    assign htif.io_scr_rdata_6 = {2{$random}};
    assign htif.io_scr_rdata_5 = {2{$random}};
    assign htif.io_scr_rdata_4 = {2{$random}};
    assign htif.io_scr_rdata_3 = {2{$random}};
    assign htif.io_scr_rdata_2 = {2{$random}};
  `endif
  FPGAOuterMemorySystem outmemsys(.clk(clk), .reset(reset),
       .io_tiles_0_acquire_ready( outmemsys_io_tiles_0_acquire_ready ),
       .io_tiles_0_acquire_valid( Queue_0_io_deq_valid ),
       .io_tiles_0_acquire_bits_header_src( Queue_0_io_deq_bits_header_src ),
       .io_tiles_0_acquire_bits_header_dst( Queue_0_io_deq_bits_header_dst ),
       .io_tiles_0_acquire_bits_payload_addr( Queue_0_io_deq_bits_payload_addr ),
       .io_tiles_0_acquire_bits_payload_client_xact_id( Queue_0_io_deq_bits_payload_client_xact_id ),
       .io_tiles_0_acquire_bits_payload_data( Queue_0_io_deq_bits_payload_data ),
       .io_tiles_0_acquire_bits_payload_a_type( Queue_0_io_deq_bits_payload_a_type ),
       .io_tiles_0_acquire_bits_payload_write_mask( Queue_0_io_deq_bits_payload_write_mask ),
       .io_tiles_0_acquire_bits_payload_subword_addr( Queue_0_io_deq_bits_payload_subword_addr ),
       .io_tiles_0_acquire_bits_payload_atomic_opcode( Queue_0_io_deq_bits_payload_atomic_opcode ),
       .io_tiles_0_grant_ready( Queue_3_io_enq_ready ),
       .io_tiles_0_grant_valid( outmemsys_io_tiles_0_grant_valid ),
       .io_tiles_0_grant_bits_header_src( outmemsys_io_tiles_0_grant_bits_header_src ),
       .io_tiles_0_grant_bits_header_dst( outmemsys_io_tiles_0_grant_bits_header_dst ),
       .io_tiles_0_grant_bits_payload_data( outmemsys_io_tiles_0_grant_bits_payload_data ),
       .io_tiles_0_grant_bits_payload_client_xact_id( outmemsys_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tiles_0_grant_bits_payload_master_xact_id( outmemsys_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_tiles_0_grant_bits_payload_g_type( outmemsys_io_tiles_0_grant_bits_payload_g_type ),
       .io_tiles_0_finish_ready( outmemsys_io_tiles_0_finish_ready ),
       .io_tiles_0_finish_valid( Queue_2_io_deq_valid ),
       .io_tiles_0_finish_bits_header_src( Queue_2_io_deq_bits_header_src ),
       .io_tiles_0_finish_bits_header_dst( Queue_2_io_deq_bits_header_dst ),
       .io_tiles_0_finish_bits_payload_master_xact_id( Queue_2_io_deq_bits_payload_master_xact_id ),
       .io_tiles_0_probe_ready( Queue_4_io_enq_ready ),
       .io_tiles_0_probe_valid( outmemsys_io_tiles_0_probe_valid ),
       .io_tiles_0_probe_bits_header_src( outmemsys_io_tiles_0_probe_bits_header_src ),
       .io_tiles_0_probe_bits_header_dst( outmemsys_io_tiles_0_probe_bits_header_dst ),
       .io_tiles_0_probe_bits_payload_addr( outmemsys_io_tiles_0_probe_bits_payload_addr ),
       .io_tiles_0_probe_bits_payload_master_xact_id( outmemsys_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_tiles_0_probe_bits_payload_p_type( outmemsys_io_tiles_0_probe_bits_payload_p_type ),
       .io_tiles_0_release_ready( outmemsys_io_tiles_0_release_ready ),
       .io_tiles_0_release_valid( Queue_1_io_deq_valid ),
       .io_tiles_0_release_bits_header_src( Queue_1_io_deq_bits_header_src ),
       .io_tiles_0_release_bits_header_dst( Queue_1_io_deq_bits_header_dst ),
       .io_tiles_0_release_bits_payload_addr( Queue_1_io_deq_bits_payload_addr ),
       .io_tiles_0_release_bits_payload_client_xact_id( Queue_1_io_deq_bits_payload_client_xact_id ),
       .io_tiles_0_release_bits_payload_master_xact_id( Queue_1_io_deq_bits_payload_master_xact_id ),
       .io_tiles_0_release_bits_payload_data( Queue_1_io_deq_bits_payload_data ),
       .io_tiles_0_release_bits_payload_r_type( Queue_1_io_deq_bits_payload_r_type ),
       .io_htif_acquire_ready( outmemsys_io_htif_acquire_ready ),
       .io_htif_acquire_valid( Queue_5_io_deq_valid ),
       .io_htif_acquire_bits_header_src( Queue_5_io_deq_bits_header_src ),
       .io_htif_acquire_bits_header_dst( Queue_5_io_deq_bits_header_dst ),
       .io_htif_acquire_bits_payload_addr( Queue_5_io_deq_bits_payload_addr ),
       .io_htif_acquire_bits_payload_client_xact_id( Queue_5_io_deq_bits_payload_client_xact_id ),
       .io_htif_acquire_bits_payload_data( Queue_5_io_deq_bits_payload_data ),
       .io_htif_acquire_bits_payload_a_type( Queue_5_io_deq_bits_payload_a_type ),
       .io_htif_acquire_bits_payload_write_mask( Queue_5_io_deq_bits_payload_write_mask ),
       .io_htif_acquire_bits_payload_subword_addr( Queue_5_io_deq_bits_payload_subword_addr ),
       .io_htif_acquire_bits_payload_atomic_opcode( Queue_5_io_deq_bits_payload_atomic_opcode ),
       .io_htif_grant_ready( Queue_8_io_enq_ready ),
       .io_htif_grant_valid( outmemsys_io_htif_grant_valid ),
       .io_htif_grant_bits_header_src( outmemsys_io_htif_grant_bits_header_src ),
       .io_htif_grant_bits_header_dst( outmemsys_io_htif_grant_bits_header_dst ),
       .io_htif_grant_bits_payload_data( outmemsys_io_htif_grant_bits_payload_data ),
       .io_htif_grant_bits_payload_client_xact_id( outmemsys_io_htif_grant_bits_payload_client_xact_id ),
       .io_htif_grant_bits_payload_master_xact_id( outmemsys_io_htif_grant_bits_payload_master_xact_id ),
       .io_htif_grant_bits_payload_g_type( outmemsys_io_htif_grant_bits_payload_g_type ),
       .io_htif_finish_ready( outmemsys_io_htif_finish_ready ),
       .io_htif_finish_valid( Queue_7_io_deq_valid ),
       .io_htif_finish_bits_header_src( Queue_7_io_deq_bits_header_src ),
       .io_htif_finish_bits_header_dst( Queue_7_io_deq_bits_header_dst ),
       .io_htif_finish_bits_payload_master_xact_id( Queue_7_io_deq_bits_payload_master_xact_id ),
       .io_htif_probe_ready( Queue_9_io_enq_ready ),
       .io_htif_probe_valid( outmemsys_io_htif_probe_valid ),
       .io_htif_probe_bits_header_src( outmemsys_io_htif_probe_bits_header_src ),
       .io_htif_probe_bits_header_dst( outmemsys_io_htif_probe_bits_header_dst ),
       .io_htif_probe_bits_payload_addr( outmemsys_io_htif_probe_bits_payload_addr ),
       .io_htif_probe_bits_payload_master_xact_id( outmemsys_io_htif_probe_bits_payload_master_xact_id ),
       .io_htif_probe_bits_payload_p_type( outmemsys_io_htif_probe_bits_payload_p_type ),
       .io_htif_release_ready( outmemsys_io_htif_release_ready ),
       .io_htif_release_valid( Queue_6_io_deq_valid ),
       .io_htif_release_bits_header_src( Queue_6_io_deq_bits_header_src ),
       .io_htif_release_bits_header_dst( Queue_6_io_deq_bits_header_dst ),
       .io_htif_release_bits_payload_addr( Queue_6_io_deq_bits_payload_addr ),
       .io_htif_release_bits_payload_client_xact_id( Queue_6_io_deq_bits_payload_client_xact_id ),
       .io_htif_release_bits_payload_master_xact_id( Queue_6_io_deq_bits_payload_master_xact_id ),
       .io_htif_release_bits_payload_data( Queue_6_io_deq_bits_payload_data ),
       .io_htif_release_bits_payload_r_type( Queue_6_io_deq_bits_payload_r_type ),
       .io_incoherent_1( 1'h1 ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( outmemsys_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( outmemsys_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( outmemsys_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( outmemsys_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( outmemsys_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( outmemsys_io_mem_req_data_bits_data ),
       .io_mem_resp_ready( outmemsys_io_mem_resp_ready ),
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag )
  );
  Queue_8 Queue_0(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_0_io_enq_ready ),
       .io_enq_valid( T43 ),
       .io_enq_bits_header_src( T42 ),
       .io_enq_bits_header_dst( T41 ),
       .io_enq_bits_payload_addr( T40 ),
       .io_enq_bits_payload_client_xact_id( T39 ),
       .io_enq_bits_payload_data( T38 ),
       .io_enq_bits_payload_a_type( T37 ),
       .io_enq_bits_payload_write_mask( T36 ),
       .io_enq_bits_payload_subword_addr( T35 ),
       .io_enq_bits_payload_atomic_opcode( T34 ),
       .io_deq_ready( outmemsys_io_tiles_0_acquire_ready ),
       .io_deq_valid( Queue_0_io_deq_valid ),
       .io_deq_bits_header_src( Queue_0_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_0_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_0_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_0_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_0_io_deq_bits_payload_data ),
       .io_deq_bits_payload_a_type( Queue_0_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_write_mask( Queue_0_io_deq_bits_payload_write_mask ),
       .io_deq_bits_payload_subword_addr( Queue_0_io_deq_bits_payload_subword_addr ),
       .io_deq_bits_payload_atomic_opcode( Queue_0_io_deq_bits_payload_atomic_opcode )
  );
  Queue_9 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( T33 ),
       .io_enq_bits_header_src( T32 ),
       .io_enq_bits_header_dst( T31 ),
       .io_enq_bits_payload_addr( T30 ),
       .io_enq_bits_payload_client_xact_id( T29 ),
       .io_enq_bits_payload_master_xact_id( T28 ),
       .io_enq_bits_payload_data( T27 ),
       .io_enq_bits_payload_r_type( T26 ),
       .io_deq_ready( outmemsys_io_tiles_0_release_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits_header_src( Queue_1_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_1_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_1_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_1_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_1_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_data( Queue_1_io_deq_bits_payload_data ),
       .io_deq_bits_payload_r_type( Queue_1_io_deq_bits_payload_r_type )
  );
  Queue_10 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( T25 ),
       .io_enq_bits_header_src( T24 ),
       .io_enq_bits_header_dst( T23 ),
       .io_enq_bits_payload_master_xact_id( T22 ),
       .io_deq_ready( outmemsys_io_tiles_0_finish_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits_header_src( Queue_2_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_2_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( Queue_2_io_deq_bits_payload_master_xact_id )
  );
  Queue_11 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( outmemsys_io_tiles_0_grant_valid ),
       .io_enq_bits_header_src( outmemsys_io_tiles_0_grant_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_tiles_0_grant_bits_header_dst ),
       .io_enq_bits_payload_data( outmemsys_io_tiles_0_grant_bits_payload_data ),
       .io_enq_bits_payload_client_xact_id( outmemsys_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_enq_bits_payload_g_type( outmemsys_io_tiles_0_grant_bits_payload_g_type ),
       .io_deq_ready( io_tiles_0_grant_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits_header_src( Queue_3_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_3_io_deq_bits_header_dst ),
       .io_deq_bits_payload_data( Queue_3_io_deq_bits_payload_data ),
       .io_deq_bits_payload_client_xact_id( Queue_3_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_3_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_g_type( Queue_3_io_deq_bits_payload_g_type )
  );
  Queue_12 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( outmemsys_io_tiles_0_probe_valid ),
       .io_enq_bits_header_src( outmemsys_io_tiles_0_probe_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_tiles_0_probe_bits_header_dst ),
       .io_enq_bits_payload_addr( outmemsys_io_tiles_0_probe_bits_payload_addr ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_enq_bits_payload_p_type( outmemsys_io_tiles_0_probe_bits_payload_p_type ),
       .io_deq_ready( io_tiles_0_probe_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_header_src( Queue_4_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_4_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_4_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_master_xact_id( Queue_4_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_p_type( Queue_4_io_deq_bits_payload_p_type )
  );
  Queue_8 Queue_5(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_5_io_enq_ready ),
       .io_enq_valid( T21 ),
       .io_enq_bits_header_src( T20 ),
       .io_enq_bits_header_dst( T19 ),
       .io_enq_bits_payload_addr( T18 ),
       .io_enq_bits_payload_client_xact_id( T17 ),
       .io_enq_bits_payload_data( T16 ),
       .io_enq_bits_payload_a_type( T15 ),
       .io_enq_bits_payload_write_mask( T14 ),
       .io_enq_bits_payload_subword_addr( T13 ),
       .io_enq_bits_payload_atomic_opcode( T12 ),
       .io_deq_ready( outmemsys_io_htif_acquire_ready ),
       .io_deq_valid( Queue_5_io_deq_valid ),
       .io_deq_bits_header_src( Queue_5_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_5_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_5_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_5_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_5_io_deq_bits_payload_data ),
       .io_deq_bits_payload_a_type( Queue_5_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_write_mask( Queue_5_io_deq_bits_payload_write_mask ),
       .io_deq_bits_payload_subword_addr( Queue_5_io_deq_bits_payload_subword_addr ),
       .io_deq_bits_payload_atomic_opcode( Queue_5_io_deq_bits_payload_atomic_opcode )
  );
  Queue_9 Queue_6(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_6_io_enq_ready ),
       .io_enq_valid( T11 ),
       .io_enq_bits_header_src( T10 ),
       .io_enq_bits_header_dst( T9 ),
       .io_enq_bits_payload_addr( T8 ),
       .io_enq_bits_payload_client_xact_id( T7 ),
       .io_enq_bits_payload_master_xact_id( T6 ),
       .io_enq_bits_payload_data( T5 ),
       .io_enq_bits_payload_r_type( T4 ),
       .io_deq_ready( outmemsys_io_htif_release_ready ),
       .io_deq_valid( Queue_6_io_deq_valid ),
       .io_deq_bits_header_src( Queue_6_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_6_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_6_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_6_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_6_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_data( Queue_6_io_deq_bits_payload_data ),
       .io_deq_bits_payload_r_type( Queue_6_io_deq_bits_payload_r_type )
  );
  Queue_10 Queue_7(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_7_io_enq_ready ),
       .io_enq_valid( T3 ),
       .io_enq_bits_header_src( T2 ),
       .io_enq_bits_header_dst( T1 ),
       .io_enq_bits_payload_master_xact_id( T0 ),
       .io_deq_ready( outmemsys_io_htif_finish_ready ),
       .io_deq_valid( Queue_7_io_deq_valid ),
       .io_deq_bits_header_src( Queue_7_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_7_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( Queue_7_io_deq_bits_payload_master_xact_id )
  );
  Queue_11 Queue_8(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_8_io_enq_ready ),
       .io_enq_valid( outmemsys_io_htif_grant_valid ),
       .io_enq_bits_header_src( outmemsys_io_htif_grant_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_htif_grant_bits_header_dst ),
       .io_enq_bits_payload_data( outmemsys_io_htif_grant_bits_payload_data ),
       .io_enq_bits_payload_client_xact_id( outmemsys_io_htif_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_htif_grant_bits_payload_master_xact_id ),
       .io_enq_bits_payload_g_type( outmemsys_io_htif_grant_bits_payload_g_type ),
       .io_deq_ready( htif_io_mem_grant_ready ),
       .io_deq_valid( Queue_8_io_deq_valid ),
       .io_deq_bits_header_src( Queue_8_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_8_io_deq_bits_header_dst ),
       .io_deq_bits_payload_data( Queue_8_io_deq_bits_payload_data ),
       .io_deq_bits_payload_client_xact_id( Queue_8_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_8_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_g_type( Queue_8_io_deq_bits_payload_g_type )
  );
  Queue_12 Queue_9(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_9_io_enq_ready ),
       .io_enq_valid( outmemsys_io_htif_probe_valid ),
       .io_enq_bits_header_src( outmemsys_io_htif_probe_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_htif_probe_bits_header_dst ),
       .io_enq_bits_payload_addr( outmemsys_io_htif_probe_bits_payload_addr ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_htif_probe_bits_payload_master_xact_id ),
       .io_enq_bits_payload_p_type( outmemsys_io_htif_probe_bits_payload_p_type ),
       .io_deq_ready( htif_io_mem_probe_ready ),
       .io_deq_valid( Queue_9_io_deq_valid ),
       .io_deq_bits_header_src( Queue_9_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_9_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_9_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_master_xact_id( Queue_9_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_p_type( Queue_9_io_deq_bits_payload_p_type )
  );
endmodule

module Queue_13(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_rw,
    input [4:0] io_enq_bits_addr,
    input [63:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_rw,
    output[4:0] io_deq_bits_addr,
    output[63:0] io_deq_bits_data
);

  wire[63:0] T0;
  wire[69:0] T1;
  wire[68:0] T2;
  wire[63:0] T3;
  wire[69:0] T4;
  reg [69:0] ram [1:0];
  wire[69:0] T5;
  wire[69:0] T6;
  wire[69:0] T7;
  wire[68:0] T8;
  wire do_enq;
  wire T9;
  wire do_flow;
  wire T10;
  reg  enq_ptr;
  wire T11;
  wire T12;
  wire T13;
  reg  deq_ptr;
  wire T14;
  wire T15;
  wire T16;
  wire do_deq;
  wire T17;
  wire T18;
  wire[4:0] T19;
  wire T20;
  wire[4:0] T21;
  wire T22;
  wire T23;
  wire empty;
  wire T24;
  reg  maybe_full;
  wire T25;
  wire T26;
  wire T27;
  wire ptr_match;
  wire T28;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {3{$random}};
    enq_ptr = {1{$random}};
    deq_ptr = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_data = T0;
  assign T0 = T1[6'h3f:1'h0];
  assign T1 = {T20, T2};
  assign T2 = {T19, T3};
  assign T3 = T4[6'h3f:1'h0];
  assign T4 = ram[deq_ptr];
  always @(posedge clk)
    if (do_enq)
      ram[enq_ptr] <= T6;
  assign T6 = T7;
  assign T7 = {io_enq_bits_rw, T8};
  assign T8 = {io_enq_bits_addr, io_enq_bits_data};
  assign do_enq = T10 & T9;
  assign T9 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T10 = io_enq_ready & io_enq_valid;
  assign T11 = reset ? 1'h0 : T12;
  assign T12 = do_enq ? T13 : enq_ptr;
  assign T13 = enq_ptr + 1'h1;
  assign T14 = reset ? 1'h0 : T15;
  assign T15 = do_deq ? T16 : deq_ptr;
  assign T16 = deq_ptr + 1'h1;
  assign do_deq = T18 & T17;
  assign T17 = do_flow ^ 1'h1;
  assign T18 = io_deq_ready & io_deq_valid;
  assign T19 = T4[7'h44:7'h40];
  assign T20 = T4[7'h45:7'h45];
  assign io_deq_bits_addr = T21;
  assign T21 = T1[7'h44:7'h40];
  assign io_deq_bits_rw = T22;
  assign T22 = T1[7'h45:7'h45];
  assign io_deq_valid = T23;
  assign T23 = empty ^ 1'h1;
  assign empty = ptr_match & T24;
  assign T24 = maybe_full ^ 1'h1;
  assign T25 = reset ? 1'h0 : T26;
  assign T26 = T27 ? do_enq : maybe_full;
  assign T27 = do_enq != do_deq;
  assign ptr_match = enq_ptr == deq_ptr;
  assign io_enq_ready = T28;
  assign T28 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      enq_ptr <= 1'h0;
    end else if(do_enq) begin
      enq_ptr <= T13;
    end
    if(reset) begin
      deq_ptr <= 1'h0;
    end else if(do_deq) begin
      deq_ptr <= T16;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T27) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_14(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [63:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[63:0] io_deq_bits
);

  wire[63:0] T0;
  reg [63:0] ram [1:0];
  wire[63:0] T1;
  wire do_enq;
  wire T2;
  wire do_flow;
  wire T3;
  reg  enq_ptr;
  wire T4;
  wire T5;
  wire T6;
  reg  deq_ptr;
  wire T7;
  wire T8;
  wire T9;
  wire do_deq;
  wire T10;
  wire T11;
  wire T12;
  wire empty;
  wire T13;
  reg  maybe_full;
  wire T14;
  wire T15;
  wire T16;
  wire ptr_match;
  wire T17;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
    enq_ptr = {1{$random}};
    deq_ptr = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits = T0;
  assign T0 = ram[deq_ptr];
  always @(posedge clk)
    if (do_enq)
      ram[enq_ptr] <= io_enq_bits;
  assign do_enq = T3 & T2;
  assign T2 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T3 = io_enq_ready & io_enq_valid;
  assign T4 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : enq_ptr;
  assign T6 = enq_ptr + 1'h1;
  assign T7 = reset ? 1'h0 : T8;
  assign T8 = do_deq ? T9 : deq_ptr;
  assign T9 = deq_ptr + 1'h1;
  assign do_deq = T11 & T10;
  assign T10 = do_flow ^ 1'h1;
  assign T11 = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T12;
  assign T12 = empty ^ 1'h1;
  assign empty = ptr_match & T13;
  assign T13 = maybe_full ^ 1'h1;
  assign T14 = reset ? 1'h0 : T15;
  assign T15 = T16 ? do_enq : maybe_full;
  assign T16 = do_enq != do_deq;
  assign ptr_match = enq_ptr == deq_ptr;
  assign io_enq_ready = T17;
  assign T17 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      enq_ptr <= 1'h0;
    end else if(do_enq) begin
      enq_ptr <= T6;
    end
    if(reset) begin
      deq_ptr <= 1'h0;
    end else if(do_deq) begin
      deq_ptr <= T9;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T16) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_15(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits
);

  wire T0;
  reg [0:0] ram [1:0];
  wire T1;
  wire do_enq;
  wire T2;
  wire do_flow;
  wire T3;
  reg  enq_ptr;
  wire T4;
  wire T5;
  wire T6;
  reg  deq_ptr;
  wire T7;
  wire T8;
  wire T9;
  wire do_deq;
  wire T10;
  wire T11;
  wire T12;
  wire empty;
  wire T13;
  reg  maybe_full;
  wire T14;
  wire T15;
  wire T16;
  wire ptr_match;
  wire T17;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    enq_ptr = {1{$random}};
    deq_ptr = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits = T0;
  assign T0 = ram[deq_ptr];
  always @(posedge clk)
    if (do_enq)
      ram[enq_ptr] <= io_enq_bits;
  assign do_enq = T3 & T2;
  assign T2 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T3 = io_enq_ready & io_enq_valid;
  assign T4 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : enq_ptr;
  assign T6 = enq_ptr + 1'h1;
  assign T7 = reset ? 1'h0 : T8;
  assign T8 = do_deq ? T9 : deq_ptr;
  assign T9 = deq_ptr + 1'h1;
  assign do_deq = T11 & T10;
  assign T10 = do_flow ^ 1'h1;
  assign T11 = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T12;
  assign T12 = empty ^ 1'h1;
  assign empty = ptr_match & T13;
  assign T13 = maybe_full ^ 1'h1;
  assign T14 = reset ? 1'h0 : T15;
  assign T15 = T16 ? do_enq : maybe_full;
  assign T16 = do_enq != do_deq;
  assign ptr_match = enq_ptr == deq_ptr;
  assign io_enq_ready = T17;
  assign T17 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      enq_ptr <= 1'h0;
    end else if(do_enq) begin
      enq_ptr <= T6;
    end
    if(reset) begin
      deq_ptr <= 1'h0;
    end else if(do_deq) begin
      deq_ptr <= T9;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T16) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module FPGATop(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    //output io_host_debug_stats_pcr
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    output io_mem_resp_ready,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
);

  wire resetSigs_0;
  wire uncore_io_htif_0_reset;
  wire Tile_io_host_ipi_rep_ready;
  wire uncore_io_htif_0_ipi_rep_bits;
  wire uncore_io_htif_0_ipi_rep_valid;
  wire uncore_io_htif_0_ipi_req_ready;
  wire Tile_io_host_ipi_req_bits;
  wire Tile_io_host_ipi_req_valid;
  wire uncore_io_htif_0_pcr_rep_ready;
  wire[63:0] Tile_io_host_pcr_rep_bits;
  wire Tile_io_host_pcr_rep_valid;
  wire Tile_io_host_pcr_req_ready;
  wire[63:0] uncore_io_htif_0_pcr_req_bits_data;
  wire[4:0] uncore_io_htif_0_pcr_req_bits_addr;
  wire uncore_io_htif_0_pcr_req_bits_rw;
  wire uncore_io_htif_0_pcr_req_valid;
  wire Queue_3_io_enq_ready;
  wire Queue_2_io_deq_bits;
  wire Queue_2_io_deq_valid;
  wire[63:0] Queue_1_io_deq_bits;
  wire Queue_1_io_deq_valid;
  wire Queue_0_io_enq_ready;
  wire[2:0] Tile_io_tilelink_release_bits_payload_r_type;
  wire[511:0] Tile_io_tilelink_release_bits_payload_data;
  wire[3:0] Tile_io_tilelink_release_bits_payload_master_xact_id;
  wire[3:0] Tile_io_tilelink_release_bits_payload_client_xact_id;
  wire[25:0] Tile_io_tilelink_release_bits_payload_addr;
  wire[1:0] Tile_io_tilelink_release_bits_header_dst;
  wire[1:0] Tile_io_tilelink_release_bits_header_src;
  wire Tile_io_tilelink_release_valid;
  wire Tile_io_tilelink_probe_ready;
  wire[3:0] Tile_io_tilelink_finish_bits_payload_master_xact_id;
  wire[1:0] Tile_io_tilelink_finish_bits_header_dst;
  wire[1:0] Tile_io_tilelink_finish_bits_header_src;
  wire Tile_io_tilelink_finish_valid;
  wire Tile_io_tilelink_grant_ready;
  wire[3:0] Tile_io_tilelink_acquire_bits_payload_atomic_opcode;
  wire[2:0] Tile_io_tilelink_acquire_bits_payload_subword_addr;
  wire[5:0] Tile_io_tilelink_acquire_bits_payload_write_mask;
  wire[2:0] Tile_io_tilelink_acquire_bits_payload_a_type;
  wire[511:0] Tile_io_tilelink_acquire_bits_payload_data;
  wire[3:0] Tile_io_tilelink_acquire_bits_payload_client_xact_id;
  wire[25:0] Tile_io_tilelink_acquire_bits_payload_addr;
  wire[1:0] Tile_io_tilelink_acquire_bits_header_dst;
  wire[1:0] Tile_io_tilelink_acquire_bits_header_src;
  wire Tile_io_tilelink_acquire_valid;
  wire Queue_3_io_deq_bits;
  wire Queue_3_io_deq_valid;
  wire Queue_2_io_enq_ready;
  wire Queue_1_io_enq_ready;
  wire[63:0] Queue_0_io_deq_bits_data;
  wire[4:0] Queue_0_io_deq_bits_addr;
  wire Queue_0_io_deq_bits_rw;
  wire Queue_0_io_deq_valid;
  reg  R0;
  reg  R1;
  wire uncore_io_tiles_0_release_ready;
  wire[1:0] uncore_io_tiles_0_probe_bits_payload_p_type;
  wire[3:0] uncore_io_tiles_0_probe_bits_payload_master_xact_id;
  wire[25:0] uncore_io_tiles_0_probe_bits_payload_addr;
  wire[1:0] uncore_io_tiles_0_probe_bits_header_dst;
  wire[1:0] uncore_io_tiles_0_probe_bits_header_src;
  wire uncore_io_tiles_0_probe_valid;
  wire uncore_io_tiles_0_finish_ready;
  wire[3:0] uncore_io_tiles_0_grant_bits_payload_g_type;
  wire[3:0] uncore_io_tiles_0_grant_bits_payload_master_xact_id;
  wire[3:0] uncore_io_tiles_0_grant_bits_payload_client_xact_id;
  wire[511:0] uncore_io_tiles_0_grant_bits_payload_data;
  wire[1:0] uncore_io_tiles_0_grant_bits_header_dst;
  wire[1:0] uncore_io_tiles_0_grant_bits_header_src;
  wire uncore_io_tiles_0_grant_valid;
  wire uncore_io_tiles_0_acquire_ready;
  wire uncore_io_mem_resp_ready;
  wire[127:0] uncore_io_mem_req_data_bits_data;
  wire uncore_io_mem_req_data_valid;
  wire uncore_io_mem_req_cmd_bits_rw;
  wire[4:0] uncore_io_mem_req_cmd_bits_tag;
  wire[25:0] uncore_io_mem_req_cmd_bits_addr;
  wire uncore_io_mem_req_cmd_valid;
  wire[15:0] uncore_io_host_out_bits;
  wire uncore_io_host_out_valid;
  wire uncore_io_host_in_ready;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R1 = {1{$random}};
  end
`endif

  assign resetSigs_0 = uncore_io_htif_0_reset;
  assign io_mem_resp_ready = uncore_io_mem_resp_ready;
  assign io_mem_req_data_bits_data = uncore_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = uncore_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = uncore_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = uncore_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = uncore_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = uncore_io_mem_req_cmd_valid;
  assign io_host_out_bits = uncore_io_host_out_bits;
  assign io_host_out_valid = uncore_io_host_out_valid;
  assign io_host_in_ready = uncore_io_host_in_ready;
  Tile Tile(.clk(clk), .reset(resetSigs_0),
       .io_tilelink_acquire_ready( uncore_io_tiles_0_acquire_ready ),
       .io_tilelink_acquire_valid( Tile_io_tilelink_acquire_valid ),
       .io_tilelink_acquire_bits_header_src( Tile_io_tilelink_acquire_bits_header_src ),
       .io_tilelink_acquire_bits_header_dst( Tile_io_tilelink_acquire_bits_header_dst ),
       .io_tilelink_acquire_bits_payload_addr( Tile_io_tilelink_acquire_bits_payload_addr ),
       .io_tilelink_acquire_bits_payload_client_xact_id( Tile_io_tilelink_acquire_bits_payload_client_xact_id ),
       .io_tilelink_acquire_bits_payload_data( Tile_io_tilelink_acquire_bits_payload_data ),
       .io_tilelink_acquire_bits_payload_a_type( Tile_io_tilelink_acquire_bits_payload_a_type ),
       .io_tilelink_acquire_bits_payload_write_mask( Tile_io_tilelink_acquire_bits_payload_write_mask ),
       .io_tilelink_acquire_bits_payload_subword_addr( Tile_io_tilelink_acquire_bits_payload_subword_addr ),
       .io_tilelink_acquire_bits_payload_atomic_opcode( Tile_io_tilelink_acquire_bits_payload_atomic_opcode ),
       .io_tilelink_grant_ready( Tile_io_tilelink_grant_ready ),
       .io_tilelink_grant_valid( uncore_io_tiles_0_grant_valid ),
       .io_tilelink_grant_bits_header_src( uncore_io_tiles_0_grant_bits_header_src ),
       .io_tilelink_grant_bits_header_dst( uncore_io_tiles_0_grant_bits_header_dst ),
       .io_tilelink_grant_bits_payload_data( uncore_io_tiles_0_grant_bits_payload_data ),
       .io_tilelink_grant_bits_payload_client_xact_id( uncore_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tilelink_grant_bits_payload_master_xact_id( uncore_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_tilelink_grant_bits_payload_g_type( uncore_io_tiles_0_grant_bits_payload_g_type ),
       .io_tilelink_finish_ready( uncore_io_tiles_0_finish_ready ),
       .io_tilelink_finish_valid( Tile_io_tilelink_finish_valid ),
       .io_tilelink_finish_bits_header_src( Tile_io_tilelink_finish_bits_header_src ),
       .io_tilelink_finish_bits_header_dst( Tile_io_tilelink_finish_bits_header_dst ),
       .io_tilelink_finish_bits_payload_master_xact_id( Tile_io_tilelink_finish_bits_payload_master_xact_id ),
       .io_tilelink_probe_ready( Tile_io_tilelink_probe_ready ),
       .io_tilelink_probe_valid( uncore_io_tiles_0_probe_valid ),
       .io_tilelink_probe_bits_header_src( uncore_io_tiles_0_probe_bits_header_src ),
       .io_tilelink_probe_bits_header_dst( uncore_io_tiles_0_probe_bits_header_dst ),
       .io_tilelink_probe_bits_payload_addr( uncore_io_tiles_0_probe_bits_payload_addr ),
       .io_tilelink_probe_bits_payload_master_xact_id( uncore_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_tilelink_probe_bits_payload_p_type( uncore_io_tiles_0_probe_bits_payload_p_type ),
       .io_tilelink_release_ready( uncore_io_tiles_0_release_ready ),
       .io_tilelink_release_valid( Tile_io_tilelink_release_valid ),
       .io_tilelink_release_bits_header_src( Tile_io_tilelink_release_bits_header_src ),
       .io_tilelink_release_bits_header_dst( Tile_io_tilelink_release_bits_header_dst ),
       .io_tilelink_release_bits_payload_addr( Tile_io_tilelink_release_bits_payload_addr ),
       .io_tilelink_release_bits_payload_client_xact_id( Tile_io_tilelink_release_bits_payload_client_xact_id ),
       .io_tilelink_release_bits_payload_master_xact_id( Tile_io_tilelink_release_bits_payload_master_xact_id ),
       .io_tilelink_release_bits_payload_data( Tile_io_tilelink_release_bits_payload_data ),
       .io_tilelink_release_bits_payload_r_type( Tile_io_tilelink_release_bits_payload_r_type ),
       .io_host_reset( R0 ),
       .io_host_id( 1'h0 ),
       .io_host_pcr_req_ready( Tile_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( Queue_0_io_deq_valid ),
       .io_host_pcr_req_bits_rw( Queue_0_io_deq_bits_rw ),
       .io_host_pcr_req_bits_addr( Queue_0_io_deq_bits_addr ),
       .io_host_pcr_req_bits_data( Queue_0_io_deq_bits_data ),
       .io_host_pcr_rep_ready( Queue_1_io_enq_ready ),
       .io_host_pcr_rep_valid( Tile_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( Tile_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( Queue_2_io_enq_ready ),
       .io_host_ipi_req_valid( Tile_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( Tile_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( Tile_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( Queue_3_io_deq_valid ),
       .io_host_ipi_rep_bits( Queue_3_io_deq_bits )
       //.io_host_debug_stats_pcr(  )
  );
  FPGAUncore uncore(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( uncore_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( uncore_io_host_out_valid ),
       .io_host_out_bits( uncore_io_host_out_bits ),
       //.io_host_debug_stats_pcr(  )
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( uncore_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( uncore_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( uncore_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( uncore_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( uncore_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( uncore_io_mem_req_data_bits_data ),
       .io_mem_resp_ready( uncore_io_mem_resp_ready ),
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag ),
       .io_tiles_0_acquire_ready( uncore_io_tiles_0_acquire_ready ),
       .io_tiles_0_acquire_valid( Tile_io_tilelink_acquire_valid ),
       .io_tiles_0_acquire_bits_header_src( Tile_io_tilelink_acquire_bits_header_src ),
       .io_tiles_0_acquire_bits_header_dst( Tile_io_tilelink_acquire_bits_header_dst ),
       .io_tiles_0_acquire_bits_payload_addr( Tile_io_tilelink_acquire_bits_payload_addr ),
       .io_tiles_0_acquire_bits_payload_client_xact_id( Tile_io_tilelink_acquire_bits_payload_client_xact_id ),
       .io_tiles_0_acquire_bits_payload_data( Tile_io_tilelink_acquire_bits_payload_data ),
       .io_tiles_0_acquire_bits_payload_a_type( Tile_io_tilelink_acquire_bits_payload_a_type ),
       .io_tiles_0_acquire_bits_payload_write_mask( Tile_io_tilelink_acquire_bits_payload_write_mask ),
       .io_tiles_0_acquire_bits_payload_subword_addr( Tile_io_tilelink_acquire_bits_payload_subword_addr ),
       .io_tiles_0_acquire_bits_payload_atomic_opcode( Tile_io_tilelink_acquire_bits_payload_atomic_opcode ),
       .io_tiles_0_grant_ready( Tile_io_tilelink_grant_ready ),
       .io_tiles_0_grant_valid( uncore_io_tiles_0_grant_valid ),
       .io_tiles_0_grant_bits_header_src( uncore_io_tiles_0_grant_bits_header_src ),
       .io_tiles_0_grant_bits_header_dst( uncore_io_tiles_0_grant_bits_header_dst ),
       .io_tiles_0_grant_bits_payload_data( uncore_io_tiles_0_grant_bits_payload_data ),
       .io_tiles_0_grant_bits_payload_client_xact_id( uncore_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tiles_0_grant_bits_payload_master_xact_id( uncore_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_tiles_0_grant_bits_payload_g_type( uncore_io_tiles_0_grant_bits_payload_g_type ),
       .io_tiles_0_finish_ready( uncore_io_tiles_0_finish_ready ),
       .io_tiles_0_finish_valid( Tile_io_tilelink_finish_valid ),
       .io_tiles_0_finish_bits_header_src( Tile_io_tilelink_finish_bits_header_src ),
       .io_tiles_0_finish_bits_header_dst( Tile_io_tilelink_finish_bits_header_dst ),
       .io_tiles_0_finish_bits_payload_master_xact_id( Tile_io_tilelink_finish_bits_payload_master_xact_id ),
       .io_tiles_0_probe_ready( Tile_io_tilelink_probe_ready ),
       .io_tiles_0_probe_valid( uncore_io_tiles_0_probe_valid ),
       .io_tiles_0_probe_bits_header_src( uncore_io_tiles_0_probe_bits_header_src ),
       .io_tiles_0_probe_bits_header_dst( uncore_io_tiles_0_probe_bits_header_dst ),
       .io_tiles_0_probe_bits_payload_addr( uncore_io_tiles_0_probe_bits_payload_addr ),
       .io_tiles_0_probe_bits_payload_master_xact_id( uncore_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_tiles_0_probe_bits_payload_p_type( uncore_io_tiles_0_probe_bits_payload_p_type ),
       .io_tiles_0_release_ready( uncore_io_tiles_0_release_ready ),
       .io_tiles_0_release_valid( Tile_io_tilelink_release_valid ),
       .io_tiles_0_release_bits_header_src( Tile_io_tilelink_release_bits_header_src ),
       .io_tiles_0_release_bits_header_dst( Tile_io_tilelink_release_bits_header_dst ),
       .io_tiles_0_release_bits_payload_addr( Tile_io_tilelink_release_bits_payload_addr ),
       .io_tiles_0_release_bits_payload_client_xact_id( Tile_io_tilelink_release_bits_payload_client_xact_id ),
       .io_tiles_0_release_bits_payload_master_xact_id( Tile_io_tilelink_release_bits_payload_master_xact_id ),
       .io_tiles_0_release_bits_payload_data( Tile_io_tilelink_release_bits_payload_data ),
       .io_tiles_0_release_bits_payload_r_type( Tile_io_tilelink_release_bits_payload_r_type ),
       .io_htif_0_reset( uncore_io_htif_0_reset ),
       //.io_htif_0_id(  )
       .io_htif_0_pcr_req_ready( Queue_0_io_enq_ready ),
       .io_htif_0_pcr_req_valid( uncore_io_htif_0_pcr_req_valid ),
       .io_htif_0_pcr_req_bits_rw( uncore_io_htif_0_pcr_req_bits_rw ),
       .io_htif_0_pcr_req_bits_addr( uncore_io_htif_0_pcr_req_bits_addr ),
       .io_htif_0_pcr_req_bits_data( uncore_io_htif_0_pcr_req_bits_data ),
       .io_htif_0_pcr_rep_ready( uncore_io_htif_0_pcr_rep_ready ),
       .io_htif_0_pcr_rep_valid( Queue_1_io_deq_valid ),
       .io_htif_0_pcr_rep_bits( Queue_1_io_deq_bits ),
       .io_htif_0_ipi_req_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_htif_0_ipi_req_valid( Queue_2_io_deq_valid ),
       .io_htif_0_ipi_req_bits( Queue_2_io_deq_bits ),
       .io_htif_0_ipi_rep_ready( Queue_3_io_enq_ready ),
       .io_htif_0_ipi_rep_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_htif_0_ipi_rep_bits( uncore_io_htif_0_ipi_rep_bits ),
       //.io_htif_0_debug_stats_pcr(  )
       .io_incoherent_0( uncore_io_htif_0_reset )
  );
  `ifndef SYNTHESIS
    assign uncore.io_htif_0_ipi_rep_bits = {1{$random}};
    assign uncore.io_htif_0_debug_stats_pcr = {1{$random}};
  `endif
  Queue_13 Queue_0(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_0_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_pcr_req_valid ),
       .io_enq_bits_rw( uncore_io_htif_0_pcr_req_bits_rw ),
       .io_enq_bits_addr( uncore_io_htif_0_pcr_req_bits_addr ),
       .io_enq_bits_data( uncore_io_htif_0_pcr_req_bits_data ),
       .io_deq_ready( Tile_io_host_pcr_req_ready ),
       .io_deq_valid( Queue_0_io_deq_valid ),
       .io_deq_bits_rw( Queue_0_io_deq_bits_rw ),
       .io_deq_bits_addr( Queue_0_io_deq_bits_addr ),
       .io_deq_bits_data( Queue_0_io_deq_bits_data )
  );
  Queue_14 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( Tile_io_host_pcr_rep_valid ),
       .io_enq_bits( Tile_io_host_pcr_rep_bits ),
       .io_deq_ready( uncore_io_htif_0_pcr_rep_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits( Queue_1_io_deq_bits )
  );
  Queue_15 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( Tile_io_host_ipi_req_valid ),
       .io_enq_bits( Tile_io_host_ipi_req_bits ),
       .io_deq_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits( Queue_2_io_deq_bits )
  );
  Queue_15 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_enq_bits( uncore_io_htif_0_ipi_rep_bits ),
       .io_deq_ready( Tile_io_host_ipi_rep_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits( Queue_3_io_deq_bits )
  );

  always @(posedge clk) begin
    R0 <= R1;
    R1 <= uncore_io_htif_0_reset;
  end
endmodule

module Queue_16(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [4:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[4:0] io_deq_bits,
    output[2:0] io_count
);

  wire[2:0] T0;
  wire[1:0] ptr_diff;
  reg [1:0] deq_ptr;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire do_deq;
  wire T4;
  wire do_flow;
  wire T5;
  reg [1:0] enq_ptr;
  wire[1:0] T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire do_enq;
  wire T9;
  wire T10;
  wire T11;
  wire ptr_match;
  reg  maybe_full;
  wire T12;
  wire T13;
  wire T14;
  wire[4:0] T15;
  reg [4:0] ram [3:0];
  wire[4:0] T16;
  wire T17;
  wire empty;
  wire T18;
  wire T19;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    deq_ptr = {1{$random}};
    enq_ptr = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T11, ptr_diff};
  assign ptr_diff = enq_ptr - deq_ptr;
  assign T1 = reset ? 2'h0 : T2;
  assign T2 = do_deq ? T3 : deq_ptr;
  assign T3 = deq_ptr + 2'h1;
  assign do_deq = T5 & T4;
  assign T4 = do_flow ^ 1'h1;
  assign do_flow = 1'h0;
  assign T5 = io_deq_ready & io_deq_valid;
  assign T6 = reset ? 2'h0 : T7;
  assign T7 = do_enq ? T8 : enq_ptr;
  assign T8 = enq_ptr + 2'h1;
  assign do_enq = T10 & T9;
  assign T9 = do_flow ^ 1'h1;
  assign T10 = io_enq_ready & io_enq_valid;
  assign T11 = maybe_full & ptr_match;
  assign ptr_match = enq_ptr == deq_ptr;
  assign T12 = reset ? 1'h0 : T13;
  assign T13 = T14 ? do_enq : maybe_full;
  assign T14 = do_enq != do_deq;
  assign io_deq_bits = T15;
  assign T15 = ram[deq_ptr];
  always @(posedge clk)
    if (do_enq)
      ram[enq_ptr] <= io_enq_bits;
  assign io_deq_valid = T17;
  assign T17 = empty ^ 1'h1;
  assign empty = ptr_match & T18;
  assign T18 = maybe_full ^ 1'h1;
  assign io_enq_ready = T19;
  assign T19 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      deq_ptr <= 2'h0;
    end else if(do_deq) begin
      deq_ptr <= T3;
    end
    if(reset) begin
      enq_ptr <= 2'h0;
    end else if(do_enq) begin
      enq_ptr <= T8;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T14) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Slave(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    input [4:0] io_addr
);

  wire T0;
  wire T1;
  reg [1:0] rf_count;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire top_io_mem_resp_ready;
  wire T6;
  wire[4:0] top_io_mem_req_cmd_bits_tag;
  wire T7;
  wire T8;
  wire top_io_mem_req_cmd_bits_rw;
  wire T9;
  wire top_io_mem_req_cmd_valid;
  wire T10;
  wire T11;
  wire[1:0] T12;
  wire[4:0] tagq_io_deq_bits;
  wire[127:0] T13;
  wire[95:0] T14;
  reg [127:0] in_reg;
  wire[127:0] T15;
  wire T16;
  wire wready_1;
  wire T17;
  wire T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  reg [1:0] in_count;
  wire[1:0] T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire[1:0] T27;
  wire T28;
  wire T29;
  reg [1:0] out_count;
  wire[1:0] T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire rvalid_2;
  wire top_io_mem_req_data_valid;
  wire T34;
  wire T35;
  wire[1:0] T36;
  wire T37;
  wire T38;
  wire[1:0] T39;
  wire T40;
  wire T41;
  wire[1:0] T42;
  wire T43;
  wire T44;
  wire[1:0] T45;
  wire[15:0] T46;
  wire T47;
  wire T48;
  wire[1:0] T49;
  wire[31:0] T50;
  wire[31:0] T51;
  wire[31:0] rdata_0;
  wire[31:0] T52;
  wire[16:0] T53;
  wire top_io_host_out_valid;
  wire[15:0] top_io_host_out_bits;
  wire[31:0] rdata_1;
  wire[31:0] T54;
  wire[27:0] T55;
  wire[1:0] T56;
  wire T57;
  wire T58;
  wire tagq_io_enq_ready;
  wire[25:0] top_io_mem_req_cmd_bits_addr;
  wire T59;
  wire[1:0] T60;
  wire[1:0] T61;
  wire[31:0] T62;
  wire[31:0] rdata_2;
  wire[31:0] T63;
  wire[127:0] T64;
  wire[7:0] T65;
  wire[127:0] top_io_mem_req_data_bits_data;
  wire[31:0] rdata_3;
  wire[31:0] T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire rvalid_0;
  wire rvalid_1;
  wire T72;
  wire[1:0] T73;
  wire[1:0] T74;
  wire T75;
  wire rvalid_3;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire wready_0;
  wire top_io_host_in_ready;
  wire T80;
  wire[1:0] T81;
  wire[1:0] T82;
  wire T83;
  wire wready_2;
  wire wready_3;
  wire T84;
  wire T85;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    rf_count = {1{$random}};
    in_reg = {4{$random}};
    in_count = {1{$random}};
    out_count = {1{$random}};
  end
`endif

  assign T0 = T6 & T1;
  assign T1 = rf_count == 2'h3;
  assign T2 = reset ? 2'h0 : T3;
  assign T3 = T5 ? T4 : rf_count;
  assign T4 = rf_count + 2'h1;
  assign T5 = top_io_mem_resp_ready & T20;
  assign T6 = top_io_mem_resp_ready & T20;
  assign T7 = T9 & T8;
  assign T8 = top_io_mem_req_cmd_bits_rw ^ 1'h1;
  assign T9 = T10 & top_io_mem_req_cmd_valid;
  assign T10 = io_out_ready & T11;
  assign T11 = T12 == 2'h1;
  assign T12 = io_addr[1'h1:1'h0];
  assign T13 = {io_in_bits, T14};
  assign T14 = in_reg[7'h7f:6'h20];
  assign T15 = T16 ? T13 : in_reg;
  assign T16 = T17 & wready_1;
  assign wready_1 = top_io_mem_resp_ready;
  assign T17 = io_in_valid & T18;
  assign T18 = T19 == 2'h1;
  assign T19 = io_addr[1'h1:1'h0];
  assign T20 = T25 & T21;
  assign T21 = in_count == 2'h3;
  assign T22 = reset ? 2'h0 : T23;
  assign T23 = T16 ? T24 : in_count;
  assign T24 = in_count + 2'h1;
  assign T25 = io_in_valid & T26;
  assign T26 = T27 == 2'h1;
  assign T27 = io_addr[1'h1:1'h0];
  assign T28 = T37 & T29;
  assign T29 = out_count == 2'h3;
  assign T30 = reset ? 2'h0 : T31;
  assign T31 = T33 ? T32 : out_count;
  assign T32 = out_count + 2'h1;
  assign T33 = T34 & rvalid_2;
  assign rvalid_2 = top_io_mem_req_data_valid;
  assign T34 = io_out_ready & T35;
  assign T35 = T36 == 2'h2;
  assign T36 = io_addr[1'h1:1'h0];
  assign T37 = io_out_ready & T38;
  assign T38 = T39 == 2'h2;
  assign T39 = io_addr[1'h1:1'h0];
  assign T40 = io_out_ready & T41;
  assign T41 = T42 == 2'h1;
  assign T42 = io_addr[1'h1:1'h0];
  assign T43 = io_out_ready & T44;
  assign T44 = T45 == 2'h0;
  assign T45 = io_addr[1'h1:1'h0];
  assign T46 = io_in_bits[4'hf:1'h0];
  assign T47 = io_in_valid & T48;
  assign T48 = T49 == 2'h0;
  assign T49 = io_addr[1'h1:1'h0];
  assign io_out_bits = T50;
  assign T50 = T69 ? T62 : T51;
  assign T51 = T59 ? rdata_1 : rdata_0;
  assign rdata_0 = T52;
  assign T52 = {15'h0, T53};
  assign T53 = {top_io_host_out_bits, top_io_host_out_valid};
  assign rdata_1 = T54;
  assign T54 = {4'h0, T55};
  assign T55 = {top_io_mem_req_cmd_bits_addr, T56};
  assign T56 = {top_io_mem_req_cmd_bits_rw, T57};
  assign T57 = top_io_mem_req_cmd_valid & T58;
  assign T58 = tagq_io_enq_ready | top_io_mem_req_cmd_bits_rw;
  assign T59 = T60[1'h0:1'h0];
  assign T60 = T61;
  assign T61 = io_addr[1'h1:1'h0];
  assign T62 = T68 ? rdata_3 : rdata_2;
  assign rdata_2 = T63;
  assign T63 = T64[5'h1f:1'h0];
  assign T64 = top_io_mem_req_data_bits_data >> T65;
  assign T65 = out_count * 6'h20;
  assign rdata_3 = T66;
  assign T66 = {30'h0, T67};
  assign T67 = {top_io_mem_req_cmd_valid, tagq_io_enq_ready};
  assign T68 = T60[1'h0:1'h0];
  assign T69 = T60[1'h1:1'h1];
  assign io_out_valid = T70;
  assign T70 = T77 ? T75 : T71;
  assign T71 = T72 ? rvalid_1 : rvalid_0;
  assign rvalid_0 = 1'h1;
  assign rvalid_1 = 1'h1;
  assign T72 = T73[1'h0:1'h0];
  assign T73 = T74;
  assign T74 = io_addr[1'h1:1'h0];
  assign T75 = T76 ? rvalid_3 : rvalid_2;
  assign rvalid_3 = 1'h1;
  assign T76 = T73[1'h0:1'h0];
  assign T77 = T73[1'h1:1'h1];
  assign io_in_ready = T78;
  assign T78 = T85 ? T83 : T79;
  assign T79 = T80 ? wready_1 : wready_0;
  assign wready_0 = top_io_host_in_ready;
  assign T80 = T81[1'h0:1'h0];
  assign T81 = T82;
  assign T82 = io_addr[1'h1:1'h0];
  assign T83 = T84 ? wready_3 : wready_2;
  assign wready_2 = 1'h1;
  assign wready_3 = 1'h1;
  assign T84 = T81[1'h0:1'h0];
  assign T85 = T81[1'h1:1'h1];
  FPGATop top(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( top_io_host_in_ready ),
       .io_host_in_valid( T47 ),
       .io_host_in_bits( T46 ),
       .io_host_out_ready( T43 ),
       .io_host_out_valid( top_io_host_out_valid ),
       .io_host_out_bits( top_io_host_out_bits ),
       //.io_host_debug_stats_pcr(  )
       .io_mem_req_cmd_ready( T40 ),
       .io_mem_req_cmd_valid( top_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( top_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( top_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( top_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( T28 ),
       .io_mem_req_data_valid( top_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( top_io_mem_req_data_bits_data ),
       .io_mem_resp_ready( top_io_mem_resp_ready ),
       .io_mem_resp_valid( T20 ),
       .io_mem_resp_bits_data( T13 ),
       .io_mem_resp_bits_tag( tagq_io_deq_bits )
  );
  Queue_16 tagq(.clk(clk), .reset(reset),
       .io_enq_ready( tagq_io_enq_ready ),
       .io_enq_valid( T7 ),
       .io_enq_bits( top_io_mem_req_cmd_bits_tag ),
       .io_deq_ready( T0 ),
       //.io_deq_valid(  )
       .io_deq_bits( tagq_io_deq_bits )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      rf_count <= 2'h0;
    end else if(T5) begin
      rf_count <= T4;
    end
    if(T16) begin
      in_reg <= T13;
    end
    if(reset) begin
      in_count <= 2'h0;
    end else if(T16) begin
      in_count <= T24;
    end
    if(reset) begin
      out_count <= 2'h0;
    end else if(T33) begin
      out_count <= T32;
    end
  end
endmodule

